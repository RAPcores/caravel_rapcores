magic
tech sky130A
magscale 1 2
timestamp 1607962800
<< locali >>
rect 154313 676243 154347 685797
rect 218989 666587 219023 676141
rect 219265 647275 219299 656829
rect 219357 616879 219391 626501
rect 219081 608719 219115 611405
rect 219265 601579 219299 608549
rect 219173 589339 219207 598893
rect 154313 579751 154347 589237
rect 364349 579683 364383 589237
rect 218897 569959 218931 579581
rect 364441 563091 364475 569857
rect 218897 550647 218931 553401
rect 154405 521679 154439 531233
rect 154405 502367 154439 511921
rect 218897 396083 218931 405637
rect 218805 354807 218839 360213
rect 359289 360111 359323 365653
rect 218989 350455 219023 354637
rect 358829 251243 358863 260797
rect 358921 234651 358955 241417
<< viali >>
rect 154313 685797 154347 685831
rect 154313 676209 154347 676243
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 219357 626501 219391 626535
rect 219357 616845 219391 616879
rect 219081 611405 219115 611439
rect 219081 608685 219115 608719
rect 219265 608549 219299 608583
rect 219265 601545 219299 601579
rect 219173 598893 219207 598927
rect 219173 589305 219207 589339
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 364349 589237 364383 589271
rect 364349 579649 364383 579683
rect 218897 579581 218931 579615
rect 218897 569925 218931 569959
rect 364441 569857 364475 569891
rect 364441 563057 364475 563091
rect 218897 553401 218931 553435
rect 218897 550613 218931 550647
rect 154405 531233 154439 531267
rect 154405 521645 154439 521679
rect 154405 511921 154439 511955
rect 154405 502333 154439 502367
rect 218897 405637 218931 405671
rect 218897 396049 218931 396083
rect 359289 365653 359323 365687
rect 218805 360213 218839 360247
rect 359289 360077 359323 360111
rect 218805 354773 218839 354807
rect 218989 354637 219023 354671
rect 218989 350421 219023 350455
rect 358829 260797 358863 260831
rect 358829 251209 358863 251243
rect 358921 241417 358955 241451
rect 358921 234617 358955 234651
<< metal1 >>
rect 295242 700544 295248 700596
rect 295300 700584 295306 700596
rect 348786 700584 348792 700596
rect 295300 700556 348792 700584
rect 295300 700544 295306 700556
rect 348786 700544 348792 700556
rect 348844 700544 348850 700596
rect 229002 700476 229008 700528
rect 229060 700516 229066 700528
rect 300118 700516 300124 700528
rect 229060 700488 300124 700516
rect 229060 700476 229066 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 283834 700408 283840 700460
rect 283892 700448 283898 700460
rect 358906 700448 358912 700460
rect 283892 700420 358912 700448
rect 283892 700408 283898 700420
rect 358906 700408 358912 700420
rect 358964 700408 358970 700460
rect 366358 700408 366364 700460
rect 366416 700448 366422 700460
rect 413646 700448 413652 700460
rect 366416 700420 413652 700448
rect 366416 700408 366422 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 240042 700340 240048 700392
rect 240100 700380 240106 700392
rect 543458 700380 543464 700392
rect 240100 700352 543464 700380
rect 240100 700340 240106 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 358814 700312 358820 700324
rect 24360 700284 358820 700312
rect 24360 700272 24366 700284
rect 358814 700272 358820 700284
rect 358872 700272 358878 700324
rect 363598 700272 363604 700324
rect 363656 700312 363662 700324
rect 478506 700312 478512 700324
rect 363656 700284 478512 700312
rect 363656 700272 363662 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 218974 694152 218980 694204
rect 219032 694192 219038 694204
rect 219158 694192 219164 694204
rect 219032 694164 219164 694192
rect 219032 694152 219038 694164
rect 219158 694152 219164 694164
rect 219216 694152 219222 694204
rect 364334 692792 364340 692844
rect 364392 692832 364398 692844
rect 365070 692832 365076 692844
rect 364392 692804 365076 692832
rect 364392 692792 364398 692804
rect 365070 692792 365076 692804
rect 365128 692792 365134 692844
rect 219158 688684 219164 688696
rect 219084 688656 219164 688684
rect 219084 688628 219112 688656
rect 219158 688644 219164 688656
rect 219216 688644 219222 688696
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 219066 688576 219072 688628
rect 219124 688576 219130 688628
rect 362218 685856 362224 685908
rect 362276 685896 362282 685908
rect 580166 685896 580172 685908
rect 362276 685868 580172 685896
rect 362276 685856 362282 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 364334 673480 364340 673532
rect 364392 673520 364398 673532
rect 364518 673520 364524 673532
rect 364392 673492 364524 673520
rect 364392 673480 364398 673492
rect 364518 673480 364524 673492
rect 364576 673480 364582 673532
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 364334 634788 364340 634840
rect 364392 634828 364398 634840
rect 364518 634828 364524 634840
rect 364392 634800 364524 634828
rect 364392 634788 364398 634800
rect 364518 634788 364524 634800
rect 364576 634788 364582 634840
rect 219342 626532 219348 626544
rect 219303 626504 219348 626532
rect 219342 626492 219348 626504
rect 219400 626492 219406 626544
rect 219342 616876 219348 616888
rect 219303 616848 219348 616876
rect 219342 616836 219348 616848
rect 219400 616836 219406 616888
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 364334 615476 364340 615528
rect 364392 615516 364398 615528
rect 364518 615516 364524 615528
rect 364392 615488 364524 615516
rect 364392 615476 364398 615488
rect 364518 615476 364524 615488
rect 364576 615476 364582 615528
rect 219069 611439 219127 611445
rect 219069 611405 219081 611439
rect 219115 611436 219127 611439
rect 219342 611436 219348 611448
rect 219115 611408 219348 611436
rect 219115 611405 219127 611408
rect 219069 611399 219127 611405
rect 219342 611396 219348 611408
rect 219400 611396 219406 611448
rect 219066 608716 219072 608728
rect 219027 608688 219072 608716
rect 219066 608676 219072 608688
rect 219124 608676 219130 608728
rect 219066 608540 219072 608592
rect 219124 608580 219130 608592
rect 219253 608583 219311 608589
rect 219253 608580 219265 608583
rect 219124 608552 219265 608580
rect 219124 608540 219130 608552
rect 219253 608549 219265 608552
rect 219299 608549 219311 608583
rect 219253 608543 219311 608549
rect 219250 601576 219256 601588
rect 219211 601548 219256 601576
rect 219250 601536 219256 601548
rect 219308 601536 219314 601588
rect 219161 598927 219219 598933
rect 219161 598893 219173 598927
rect 219207 598924 219219 598927
rect 219250 598924 219256 598936
rect 219207 598896 219256 598924
rect 219207 598893 219219 598896
rect 219161 598887 219219 598893
rect 219250 598884 219256 598896
rect 219308 598884 219314 598936
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 364334 596164 364340 596216
rect 364392 596204 364398 596216
rect 364518 596204 364524 596216
rect 364392 596176 364524 596204
rect 364392 596164 364398 596176
rect 364518 596164 364524 596176
rect 364576 596164 364582 596216
rect 362310 592016 362316 592068
rect 362368 592056 362374 592068
rect 580166 592056 580172 592068
rect 362368 592028 580172 592056
rect 362368 592016 362374 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 219158 589336 219164 589348
rect 219119 589308 219164 589336
rect 219158 589296 219164 589308
rect 219216 589296 219222 589348
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 364337 589271 364395 589277
rect 364337 589237 364349 589271
rect 364383 589268 364395 589271
rect 364426 589268 364432 589280
rect 364383 589240 364432 589268
rect 364383 589237 364395 589240
rect 364337 589231 364395 589237
rect 364426 589228 364432 589240
rect 364484 589228 364490 589280
rect 218974 582360 218980 582412
rect 219032 582400 219038 582412
rect 219158 582400 219164 582412
rect 219032 582372 219164 582400
rect 219032 582360 219038 582372
rect 219158 582360 219164 582372
rect 219216 582360 219222 582412
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 364334 579680 364340 579692
rect 364295 579652 364340 579680
rect 364334 579640 364340 579652
rect 364392 579640 364398 579692
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 218885 579615 218943 579621
rect 218885 579581 218897 579615
rect 218931 579612 218943 579615
rect 218974 579612 218980 579624
rect 218931 579584 218980 579612
rect 218931 579581 218943 579584
rect 218885 579575 218943 579581
rect 218974 579572 218980 579584
rect 219032 579572 219038 579624
rect 218882 569956 218888 569968
rect 218843 569928 218888 569956
rect 218882 569916 218888 569928
rect 218940 569916 218946 569968
rect 364426 569888 364432 569900
rect 364387 569860 364432 569888
rect 364426 569848 364432 569860
rect 364484 569848 364490 569900
rect 3326 567196 3332 567248
rect 3384 567236 3390 567248
rect 358998 567236 359004 567248
rect 3384 567208 359004 567236
rect 3384 567196 3390 567208
rect 358998 567196 359004 567208
rect 359056 567196 359062 567248
rect 218882 563048 218888 563100
rect 218940 563048 218946 563100
rect 364429 563091 364487 563097
rect 364429 563057 364441 563091
rect 364475 563088 364487 563091
rect 364610 563088 364616 563100
rect 364475 563060 364616 563088
rect 364475 563057 364487 563060
rect 364429 563051 364487 563057
rect 364610 563048 364616 563060
rect 364668 563048 364674 563100
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 218900 562952 218928 563048
rect 218974 562952 218980 562964
rect 218900 562924 218980 562952
rect 218974 562912 218980 562924
rect 219032 562912 219038 562964
rect 218882 553432 218888 553444
rect 218843 553404 218888 553432
rect 218882 553392 218888 553404
rect 218940 553392 218946 553444
rect 218882 550644 218888 550656
rect 218843 550616 218888 550644
rect 218882 550604 218888 550616
rect 218940 550604 218946 550656
rect 364426 550604 364432 550656
rect 364484 550644 364490 550656
rect 364702 550644 364708 550656
rect 364484 550616 364708 550644
rect 364484 550604 364490 550616
rect 364702 550604 364708 550616
rect 364760 550604 364766 550656
rect 362402 545096 362408 545148
rect 362460 545136 362466 545148
rect 580166 545136 580172 545148
rect 362460 545108 580172 545136
rect 362460 545096 362466 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 364702 543844 364708 543856
rect 364628 543816 364708 543844
rect 218882 543736 218888 543788
rect 218940 543736 218946 543788
rect 218900 543640 218928 543736
rect 364628 543720 364656 543816
rect 364702 543804 364708 543816
rect 364760 543804 364766 543856
rect 364610 543668 364616 543720
rect 364668 543668 364674 543720
rect 218974 543640 218980 543652
rect 218900 543612 218980 543640
rect 218974 543600 218980 543612
rect 219032 543600 219038 543652
rect 364426 531292 364432 531344
rect 364484 531332 364490 531344
rect 364702 531332 364708 531344
rect 364484 531304 364708 531332
rect 364484 531292 364490 531304
rect 364702 531292 364708 531304
rect 364760 531292 364766 531344
rect 154390 531264 154396 531276
rect 154351 531236 154396 531264
rect 154390 531224 154396 531236
rect 154448 531224 154454 531276
rect 364702 524532 364708 524544
rect 364628 524504 364708 524532
rect 364628 524408 364656 524504
rect 364702 524492 364708 524504
rect 364760 524492 364766 524544
rect 364610 524356 364616 524408
rect 364668 524356 364674 524408
rect 218974 524288 218980 524340
rect 219032 524328 219038 524340
rect 219158 524328 219164 524340
rect 219032 524300 219164 524328
rect 219032 524288 219038 524300
rect 219158 524288 219164 524300
rect 219216 524288 219222 524340
rect 154393 521679 154451 521685
rect 154393 521645 154405 521679
rect 154439 521676 154451 521679
rect 154482 521676 154488 521688
rect 154439 521648 154488 521676
rect 154439 521645 154451 521648
rect 154393 521639 154451 521645
rect 154482 521636 154488 521648
rect 154540 521636 154546 521688
rect 364426 511980 364432 512032
rect 364484 512020 364490 512032
rect 364702 512020 364708 512032
rect 364484 511992 364708 512020
rect 364484 511980 364490 511992
rect 364702 511980 364708 511992
rect 364760 511980 364766 512032
rect 154390 511952 154396 511964
rect 154351 511924 154396 511952
rect 154390 511912 154396 511924
rect 154448 511912 154454 511964
rect 154393 502367 154451 502373
rect 154393 502333 154405 502367
rect 154439 502364 154451 502367
rect 154482 502364 154488 502376
rect 154439 502336 154488 502364
rect 154439 502333 154451 502336
rect 154393 502327 154451 502333
rect 154482 502324 154488 502336
rect 154540 502324 154546 502376
rect 218882 502324 218888 502376
rect 218940 502364 218946 502376
rect 219342 502364 219348 502376
rect 218940 502336 219348 502364
rect 218940 502324 218946 502336
rect 219342 502324 219348 502336
rect 219400 502324 219406 502376
rect 364518 502324 364524 502376
rect 364576 502364 364582 502376
rect 364702 502364 364708 502376
rect 364576 502336 364708 502364
rect 364576 502324 364582 502336
rect 364702 502324 364708 502336
rect 364760 502324 364766 502376
rect 3326 495456 3332 495508
rect 3384 495496 3390 495508
rect 359090 495496 359096 495508
rect 3384 495468 359096 495496
rect 3384 495456 3390 495468
rect 359090 495456 359096 495468
rect 359148 495456 359154 495508
rect 154298 485800 154304 485852
rect 154356 485800 154362 485852
rect 314562 485800 314568 485852
rect 314620 485840 314626 485852
rect 580166 485840 580172 485852
rect 314620 485812 580172 485840
rect 314620 485800 314626 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 154316 485704 154344 485800
rect 154390 485704 154396 485716
rect 154316 485676 154396 485704
rect 154390 485664 154396 485676
rect 154448 485664 154454 485716
rect 154114 482944 154120 482996
rect 154172 482984 154178 482996
rect 154390 482984 154396 482996
rect 154172 482956 154396 482984
rect 154172 482944 154178 482956
rect 154390 482944 154396 482956
rect 154448 482944 154454 482996
rect 219158 480224 219164 480276
rect 219216 480264 219222 480276
rect 219342 480264 219348 480276
rect 219216 480236 219348 480264
rect 219216 480224 219222 480236
rect 219342 480224 219348 480236
rect 219400 480224 219406 480276
rect 364334 480224 364340 480276
rect 364392 480264 364398 480276
rect 364518 480264 364524 480276
rect 364392 480236 364524 480264
rect 364392 480224 364398 480236
rect 364518 480224 364524 480236
rect 364576 480224 364582 480276
rect 313642 472676 313648 472728
rect 313700 472716 313706 472728
rect 314562 472716 314568 472728
rect 313700 472688 314568 472716
rect 313700 472676 313706 472688
rect 314562 472676 314568 472688
rect 314620 472676 314626 472728
rect 154298 472608 154304 472660
rect 154356 472648 154362 472660
rect 276474 472648 276480 472660
rect 154356 472620 276480 472648
rect 154356 472608 154362 472620
rect 276474 472608 276480 472620
rect 276532 472608 276538 472660
rect 3602 472064 3608 472116
rect 3660 472104 3666 472116
rect 257890 472104 257896 472116
rect 3660 472076 257896 472104
rect 3660 472064 3666 472076
rect 257890 472064 257896 472076
rect 257948 472064 257954 472116
rect 3694 471996 3700 472048
rect 3752 472036 3758 472048
rect 350810 472036 350816 472048
rect 3752 472008 350816 472036
rect 3752 471996 3758 472008
rect 350810 471996 350816 472008
rect 350868 471996 350874 472048
rect 219158 460912 219164 460964
rect 219216 460952 219222 460964
rect 219342 460952 219348 460964
rect 219216 460924 219348 460952
rect 219216 460912 219222 460924
rect 219342 460912 219348 460924
rect 219400 460912 219406 460964
rect 364334 460912 364340 460964
rect 364392 460952 364398 460964
rect 364518 460952 364524 460964
rect 364392 460924 364524 460952
rect 364392 460912 364398 460924
rect 364518 460912 364524 460924
rect 364576 460912 364582 460964
rect 219250 444320 219256 444372
rect 219308 444360 219314 444372
rect 219434 444360 219440 444372
rect 219308 444332 219440 444360
rect 219308 444320 219314 444332
rect 219434 444320 219440 444332
rect 219492 444320 219498 444372
rect 364334 441600 364340 441652
rect 364392 441640 364398 441652
rect 364518 441640 364524 441652
rect 364392 441612 364524 441640
rect 364392 441600 364398 441612
rect 364518 441600 364524 441612
rect 364576 441600 364582 441652
rect 359458 438880 359464 438932
rect 359516 438920 359522 438932
rect 580166 438920 580172 438932
rect 359516 438892 580172 438920
rect 359516 438880 359522 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 218974 427796 218980 427848
rect 219032 427836 219038 427848
rect 219158 427836 219164 427848
rect 219032 427808 219164 427836
rect 219032 427796 219038 427808
rect 219158 427796 219164 427808
rect 219216 427796 219222 427848
rect 218698 425008 218704 425060
rect 218756 425048 218762 425060
rect 218974 425048 218980 425060
rect 218756 425020 218980 425048
rect 218756 425008 218762 425020
rect 218974 425008 218980 425020
rect 219032 425008 219038 425060
rect 364334 422288 364340 422340
rect 364392 422328 364398 422340
rect 364518 422328 364524 422340
rect 364392 422300 364524 422328
rect 364392 422288 364398 422300
rect 364518 422288 364524 422300
rect 364576 422288 364582 422340
rect 359182 419296 359188 419348
rect 359240 419336 359246 419348
rect 359550 419336 359556 419348
rect 359240 419308 359556 419336
rect 359240 419296 359246 419308
rect 359550 419296 359556 419308
rect 359608 419296 359614 419348
rect 218882 408484 218888 408536
rect 218940 408484 218946 408536
rect 218900 408388 218928 408484
rect 218974 408388 218980 408400
rect 218900 408360 218980 408388
rect 218974 408348 218980 408360
rect 219032 408348 219038 408400
rect 218885 405671 218943 405677
rect 218885 405637 218897 405671
rect 218931 405668 218943 405671
rect 218974 405668 218980 405680
rect 218931 405640 218980 405668
rect 218931 405637 218943 405640
rect 218885 405631 218943 405637
rect 218974 405628 218980 405640
rect 219032 405628 219038 405680
rect 359182 405560 359188 405612
rect 359240 405600 359246 405612
rect 359550 405600 359556 405612
rect 359240 405572 359556 405600
rect 359240 405560 359246 405572
rect 359550 405560 359556 405572
rect 359608 405560 359614 405612
rect 364334 402976 364340 403028
rect 364392 403016 364398 403028
rect 364518 403016 364524 403028
rect 364392 402988 364524 403016
rect 364392 402976 364398 402988
rect 364518 402976 364524 402988
rect 364576 402976 364582 403028
rect 218882 396080 218888 396092
rect 218843 396052 218888 396080
rect 218882 396040 218888 396052
rect 218940 396040 218946 396092
rect 3326 395972 3332 396024
rect 3384 396012 3390 396024
rect 228358 396012 228364 396024
rect 3384 395984 217364 396012
rect 3384 395972 3390 395984
rect 217336 395944 217364 395984
rect 218992 395984 228364 396012
rect 218992 395944 219020 395984
rect 228358 395972 228364 395984
rect 228416 395972 228422 396024
rect 217336 395916 219020 395944
rect 359182 389444 359188 389496
rect 359240 389484 359246 389496
rect 359550 389484 359556 389496
rect 359240 389456 359556 389484
rect 359240 389444 359246 389456
rect 359550 389444 359556 389456
rect 359608 389444 359614 389496
rect 364334 383664 364340 383716
rect 364392 383704 364398 383716
rect 364518 383704 364524 383716
rect 364392 383676 364524 383704
rect 364392 383664 364398 383676
rect 364518 383664 364524 383676
rect 364576 383664 364582 383716
rect 359274 375368 359280 375420
rect 359332 375408 359338 375420
rect 359550 375408 359556 375420
rect 359332 375380 359556 375408
rect 359332 375368 359338 375380
rect 359550 375368 359556 375380
rect 359608 375368 359614 375420
rect 218974 372580 218980 372632
rect 219032 372620 219038 372632
rect 219158 372620 219164 372632
rect 219032 372592 219164 372620
rect 219032 372580 219038 372592
rect 219158 372580 219164 372592
rect 219216 372580 219222 372632
rect 218974 367752 218980 367804
rect 219032 367792 219038 367804
rect 219158 367792 219164 367804
rect 219032 367764 219164 367792
rect 219032 367752 219038 367764
rect 219158 367752 219164 367764
rect 219216 367752 219222 367804
rect 359274 365684 359280 365696
rect 359235 365656 359280 365684
rect 359274 365644 359280 365656
rect 359332 365644 359338 365696
rect 364334 364352 364340 364404
rect 364392 364392 364398 364404
rect 364518 364392 364524 364404
rect 364392 364364 364524 364392
rect 364392 364352 364398 364364
rect 364518 364352 364524 364364
rect 364576 364352 364582 364404
rect 218793 360247 218851 360253
rect 218793 360213 218805 360247
rect 218839 360244 218851 360247
rect 218974 360244 218980 360256
rect 218839 360216 218980 360244
rect 218839 360213 218851 360216
rect 218793 360207 218851 360213
rect 218974 360204 218980 360216
rect 219032 360204 219038 360256
rect 359182 360068 359188 360120
rect 359240 360108 359246 360120
rect 359277 360111 359335 360117
rect 359277 360108 359289 360111
rect 359240 360080 359289 360108
rect 359240 360068 359246 360080
rect 359277 360077 359289 360080
rect 359323 360077 359335 360111
rect 359277 360071 359335 360077
rect 218790 354804 218796 354816
rect 218751 354776 218796 354804
rect 218790 354764 218796 354776
rect 218848 354764 218854 354816
rect 218790 354628 218796 354680
rect 218848 354668 218854 354680
rect 218977 354671 219035 354677
rect 218977 354668 218989 354671
rect 218848 354640 218989 354668
rect 218848 354628 218854 354640
rect 218977 354637 218989 354640
rect 219023 354637 219035 354671
rect 218977 354631 219035 354637
rect 218974 350452 218980 350464
rect 218935 350424 218980 350452
rect 218974 350412 218980 350424
rect 219032 350412 219038 350464
rect 364334 345040 364340 345092
rect 364392 345080 364398 345092
rect 364518 345080 364524 345092
rect 364392 345052 364524 345080
rect 364392 345040 364398 345052
rect 364518 345040 364524 345052
rect 364576 345040 364582 345092
rect 218974 340932 218980 340944
rect 218900 340904 218980 340932
rect 218900 340876 218928 340904
rect 218974 340892 218980 340904
rect 219032 340892 219038 340944
rect 218882 340824 218888 340876
rect 218940 340824 218946 340876
rect 3510 338036 3516 338088
rect 3568 338076 3574 338088
rect 352006 338076 352012 338088
rect 3568 338048 352012 338076
rect 3568 338036 3574 338048
rect 352006 338036 352012 338048
rect 352064 338036 352070 338088
rect 3418 337968 3424 338020
rect 3476 338008 3482 338020
rect 270770 338008 270776 338020
rect 3476 337980 270776 338008
rect 3476 337968 3482 337980
rect 270770 337968 270776 337980
rect 270828 337968 270834 338020
rect 286962 337968 286968 338020
rect 287020 338008 287026 338020
rect 363598 338008 363604 338020
rect 287020 337980 363604 338008
rect 287020 337968 287026 337980
rect 363598 337968 363604 337980
rect 363656 337968 363662 338020
rect 238294 337900 238300 337952
rect 238352 337940 238358 337952
rect 359458 337940 359464 337952
rect 238352 337912 359464 337940
rect 238352 337900 238358 337912
rect 359458 337900 359464 337912
rect 359516 337900 359522 337952
rect 254486 337832 254492 337884
rect 254544 337872 254550 337884
rect 364334 337872 364340 337884
rect 254544 337844 364340 337872
rect 254544 337832 254550 337844
rect 364334 337832 364340 337844
rect 364392 337832 364398 337884
rect 218882 337764 218888 337816
rect 218940 337804 218946 337816
rect 303246 337804 303252 337816
rect 218940 337776 303252 337804
rect 218940 337764 218946 337776
rect 303246 337764 303252 337776
rect 303304 337764 303310 337816
rect 319530 337764 319536 337816
rect 319588 337804 319594 337816
rect 366358 337804 366364 337816
rect 319588 337776 366364 337804
rect 319588 337764 319594 337776
rect 366358 337764 366364 337776
rect 366416 337764 366422 337816
rect 3694 337356 3700 337408
rect 3752 337396 3758 337408
rect 335722 337396 335728 337408
rect 3752 337368 335728 337396
rect 3752 337356 3758 337368
rect 335722 337356 335728 337368
rect 335780 337356 335786 337408
rect 358814 335316 358820 335368
rect 358872 335356 358878 335368
rect 359090 335356 359096 335368
rect 358872 335328 359096 335356
rect 358872 335316 358878 335328
rect 359090 335316 359096 335328
rect 359148 335316 359154 335368
rect 358814 325592 358820 325644
rect 358872 325632 358878 325644
rect 359090 325632 359096 325644
rect 358872 325604 359096 325632
rect 358872 325592 358878 325604
rect 359090 325592 359096 325604
rect 359148 325592 359154 325644
rect 358814 316004 358820 316056
rect 358872 316044 358878 316056
rect 359090 316044 359096 316056
rect 358872 316016 359096 316044
rect 358872 316004 358878 316016
rect 359090 316004 359096 316016
rect 359148 316004 359154 316056
rect 358814 306280 358820 306332
rect 358872 306320 358878 306332
rect 359090 306320 359096 306332
rect 358872 306292 359096 306320
rect 358872 306280 358878 306292
rect 359090 306280 359096 306292
rect 359148 306280 359154 306332
rect 358814 296692 358820 296744
rect 358872 296732 358878 296744
rect 359090 296732 359096 296744
rect 358872 296704 359096 296732
rect 358872 296692 358878 296704
rect 359090 296692 359096 296704
rect 359148 296692 359154 296744
rect 358814 286968 358820 287020
rect 358872 287008 358878 287020
rect 359090 287008 359096 287020
rect 358872 286980 359096 287008
rect 358872 286968 358878 286980
rect 359090 286968 359096 286980
rect 359148 286968 359154 287020
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 358906 280140 358912 280152
rect 3476 280112 358912 280140
rect 3476 280100 3482 280112
rect 358906 280100 358912 280112
rect 358964 280100 358970 280152
rect 358814 277380 358820 277432
rect 358872 277420 358878 277432
rect 359090 277420 359096 277432
rect 358872 277392 359096 277420
rect 358872 277380 358878 277392
rect 359090 277380 359096 277392
rect 359148 277380 359154 277432
rect 358814 267724 358820 267776
rect 358872 267764 358878 267776
rect 358998 267764 359004 267776
rect 358872 267736 359004 267764
rect 358872 267724 358878 267736
rect 358998 267724 359004 267736
rect 359056 267724 359062 267776
rect 358817 260831 358875 260837
rect 358817 260797 358829 260831
rect 358863 260828 358875 260831
rect 358906 260828 358912 260840
rect 358863 260800 358912 260828
rect 358863 260797 358875 260800
rect 358817 260791 358875 260797
rect 358906 260788 358912 260800
rect 358964 260788 358970 260840
rect 358814 251240 358820 251252
rect 358775 251212 358820 251240
rect 358814 251200 358820 251212
rect 358872 251200 358878 251252
rect 358906 241448 358912 241460
rect 358867 241420 358912 241448
rect 358906 241408 358912 241420
rect 358964 241408 358970 241460
rect 358909 234651 358967 234657
rect 358909 234617 358921 234651
rect 358955 234648 358967 234651
rect 359090 234648 359096 234660
rect 358955 234620 359096 234648
rect 358955 234617 358967 234620
rect 358909 234611 358967 234617
rect 359090 234608 359096 234620
rect 359148 234608 359154 234660
rect 358906 222164 358912 222216
rect 358964 222204 358970 222216
rect 359182 222204 359188 222216
rect 358964 222176 359188 222204
rect 358964 222164 358970 222176
rect 359182 222164 359188 222176
rect 359240 222164 359246 222216
rect 359182 215404 359188 215416
rect 359108 215376 359188 215404
rect 359108 215280 359136 215376
rect 359182 215364 359188 215376
rect 359240 215364 359246 215416
rect 359090 215228 359096 215280
rect 359148 215228 359154 215280
rect 358906 202852 358912 202904
rect 358964 202892 358970 202904
rect 359182 202892 359188 202904
rect 358964 202864 359188 202892
rect 358964 202852 358970 202864
rect 359182 202852 359188 202864
rect 359240 202852 359246 202904
rect 359182 196092 359188 196104
rect 359108 196064 359188 196092
rect 359108 195968 359136 196064
rect 359182 196052 359188 196064
rect 359240 196052 359246 196104
rect 359090 195916 359096 195968
rect 359148 195916 359154 195968
rect 358906 183540 358912 183592
rect 358964 183580 358970 183592
rect 359182 183580 359188 183592
rect 358964 183552 359188 183580
rect 358964 183540 358970 183552
rect 359182 183540 359188 183552
rect 359240 183540 359246 183592
rect 358998 173884 359004 173936
rect 359056 173924 359062 173936
rect 359182 173924 359188 173936
rect 359056 173896 359188 173924
rect 359056 173884 359062 173896
rect 359182 173884 359188 173896
rect 359240 173884 359246 173936
rect 358814 151784 358820 151836
rect 358872 151824 358878 151836
rect 358998 151824 359004 151836
rect 358872 151796 359004 151824
rect 358872 151784 358878 151796
rect 358998 151784 359004 151796
rect 359056 151784 359062 151836
rect 358814 132472 358820 132524
rect 358872 132512 358878 132524
rect 358998 132512 359004 132524
rect 358872 132484 359004 132512
rect 358872 132472 358878 132484
rect 358998 132472 359004 132484
rect 359056 132472 359062 132524
rect 358814 113160 358820 113212
rect 358872 113200 358878 113212
rect 358998 113200 359004 113212
rect 358872 113172 359004 113200
rect 358872 113160 358878 113172
rect 358998 113160 359004 113172
rect 359056 113160 359062 113212
rect 358814 93848 358820 93900
rect 358872 93888 358878 93900
rect 358998 93888 359004 93900
rect 358872 93860 359004 93888
rect 358872 93848 358878 93860
rect 358998 93848 359004 93860
rect 359056 93848 359062 93900
rect 358814 74536 358820 74588
rect 358872 74576 358878 74588
rect 358998 74576 359004 74588
rect 358872 74548 359004 74576
rect 358872 74536 358878 74548
rect 358998 74536 359004 74548
rect 359056 74536 359062 74588
rect 358814 55224 358820 55276
rect 358872 55264 358878 55276
rect 358998 55264 359004 55276
rect 358872 55236 359004 55264
rect 358872 55224 358878 55236
rect 358998 55224 359004 55236
rect 359056 55224 359062 55276
rect 358814 35912 358820 35964
rect 358872 35952 358878 35964
rect 358998 35952 359004 35964
rect 358872 35924 359004 35952
rect 358872 35912 358878 35924
rect 358998 35912 359004 35924
rect 359056 35912 359062 35964
rect 358814 16600 358820 16652
rect 358872 16640 358878 16652
rect 358998 16640 359004 16652
rect 358872 16612 359004 16640
rect 358872 16600 358878 16612
rect 358998 16600 359004 16612
rect 359056 16600 359062 16652
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 358998 3448 359004 3460
rect 624 3420 359004 3448
rect 624 3408 630 3420
rect 358998 3408 359004 3420
rect 359056 3408 359062 3460
<< via1 >>
rect 295248 700544 295300 700596
rect 348792 700544 348844 700596
rect 229008 700476 229060 700528
rect 300124 700476 300176 700528
rect 283840 700408 283892 700460
rect 358912 700408 358964 700460
rect 366364 700408 366416 700460
rect 413652 700408 413704 700460
rect 240048 700340 240100 700392
rect 543464 700340 543516 700392
rect 24308 700272 24360 700324
rect 358820 700272 358872 700324
rect 363604 700272 363656 700324
rect 478512 700272 478564 700324
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 218980 694152 219032 694204
rect 219164 694152 219216 694204
rect 364340 692792 364392 692844
rect 365076 692792 365128 692844
rect 219164 688644 219216 688696
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 219072 688576 219124 688628
rect 362224 685856 362276 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 364340 673480 364392 673532
rect 364524 673480 364576 673532
rect 219072 666544 219124 666596
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 219348 656820 219400 656872
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 219256 640364 219308 640416
rect 219072 640228 219124 640280
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 364340 634788 364392 634840
rect 364524 634788 364576 634840
rect 219348 626535 219400 626544
rect 219348 626501 219357 626535
rect 219357 626501 219391 626535
rect 219391 626501 219400 626535
rect 219348 626492 219400 626501
rect 219348 616879 219400 616888
rect 219348 616845 219357 616879
rect 219357 616845 219391 616879
rect 219391 616845 219400 616879
rect 219348 616836 219400 616845
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 364340 615476 364392 615528
rect 364524 615476 364576 615528
rect 219348 611396 219400 611448
rect 219072 608719 219124 608728
rect 219072 608685 219081 608719
rect 219081 608685 219115 608719
rect 219115 608685 219124 608719
rect 219072 608676 219124 608685
rect 219072 608540 219124 608592
rect 219256 601579 219308 601588
rect 219256 601545 219265 601579
rect 219265 601545 219299 601579
rect 219299 601545 219308 601579
rect 219256 601536 219308 601545
rect 219256 598884 219308 598936
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 364340 596164 364392 596216
rect 364524 596164 364576 596216
rect 362316 592016 362368 592068
rect 580172 592016 580224 592068
rect 219164 589339 219216 589348
rect 219164 589305 219173 589339
rect 219173 589305 219207 589339
rect 219207 589305 219216 589339
rect 219164 589296 219216 589305
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 364432 589228 364484 589280
rect 218980 582360 219032 582412
rect 219164 582360 219216 582412
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 364340 579683 364392 579692
rect 364340 579649 364349 579683
rect 364349 579649 364383 579683
rect 364383 579649 364392 579683
rect 364340 579640 364392 579649
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 218980 579572 219032 579624
rect 218888 569959 218940 569968
rect 218888 569925 218897 569959
rect 218897 569925 218931 569959
rect 218931 569925 218940 569959
rect 218888 569916 218940 569925
rect 364432 569891 364484 569900
rect 364432 569857 364441 569891
rect 364441 569857 364475 569891
rect 364475 569857 364484 569891
rect 364432 569848 364484 569857
rect 3332 567196 3384 567248
rect 359004 567196 359056 567248
rect 218888 563048 218940 563100
rect 364616 563048 364668 563100
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 218980 562912 219032 562964
rect 218888 553435 218940 553444
rect 218888 553401 218897 553435
rect 218897 553401 218931 553435
rect 218931 553401 218940 553435
rect 218888 553392 218940 553401
rect 218888 550647 218940 550656
rect 218888 550613 218897 550647
rect 218897 550613 218931 550647
rect 218931 550613 218940 550647
rect 218888 550604 218940 550613
rect 364432 550604 364484 550656
rect 364708 550604 364760 550656
rect 362408 545096 362460 545148
rect 580172 545096 580224 545148
rect 218888 543736 218940 543788
rect 364708 543804 364760 543856
rect 364616 543668 364668 543720
rect 218980 543600 219032 543652
rect 364432 531292 364484 531344
rect 364708 531292 364760 531344
rect 154396 531267 154448 531276
rect 154396 531233 154405 531267
rect 154405 531233 154439 531267
rect 154439 531233 154448 531267
rect 154396 531224 154448 531233
rect 364708 524492 364760 524544
rect 364616 524356 364668 524408
rect 218980 524288 219032 524340
rect 219164 524288 219216 524340
rect 154488 521636 154540 521688
rect 364432 511980 364484 512032
rect 364708 511980 364760 512032
rect 154396 511955 154448 511964
rect 154396 511921 154405 511955
rect 154405 511921 154439 511955
rect 154439 511921 154448 511955
rect 154396 511912 154448 511921
rect 154488 502324 154540 502376
rect 218888 502324 218940 502376
rect 219348 502324 219400 502376
rect 364524 502324 364576 502376
rect 364708 502324 364760 502376
rect 3332 495456 3384 495508
rect 359096 495456 359148 495508
rect 154304 485800 154356 485852
rect 314568 485800 314620 485852
rect 580172 485800 580224 485852
rect 154396 485664 154448 485716
rect 154120 482944 154172 482996
rect 154396 482944 154448 482996
rect 219164 480224 219216 480276
rect 219348 480224 219400 480276
rect 364340 480224 364392 480276
rect 364524 480224 364576 480276
rect 313648 472676 313700 472728
rect 314568 472676 314620 472728
rect 154304 472608 154356 472660
rect 276480 472608 276532 472660
rect 3608 472064 3660 472116
rect 257896 472064 257948 472116
rect 3700 471996 3752 472048
rect 350816 471996 350868 472048
rect 219164 460912 219216 460964
rect 219348 460912 219400 460964
rect 364340 460912 364392 460964
rect 364524 460912 364576 460964
rect 219256 444320 219308 444372
rect 219440 444320 219492 444372
rect 364340 441600 364392 441652
rect 364524 441600 364576 441652
rect 359464 438880 359516 438932
rect 580172 438880 580224 438932
rect 218980 427796 219032 427848
rect 219164 427796 219216 427848
rect 218704 425008 218756 425060
rect 218980 425008 219032 425060
rect 364340 422288 364392 422340
rect 364524 422288 364576 422340
rect 359188 419296 359240 419348
rect 359556 419296 359608 419348
rect 218888 408484 218940 408536
rect 218980 408348 219032 408400
rect 218980 405628 219032 405680
rect 359188 405560 359240 405612
rect 359556 405560 359608 405612
rect 364340 402976 364392 403028
rect 364524 402976 364576 403028
rect 218888 396083 218940 396092
rect 218888 396049 218897 396083
rect 218897 396049 218931 396083
rect 218931 396049 218940 396083
rect 218888 396040 218940 396049
rect 3332 395972 3384 396024
rect 228364 395972 228416 396024
rect 359188 389444 359240 389496
rect 359556 389444 359608 389496
rect 364340 383664 364392 383716
rect 364524 383664 364576 383716
rect 359280 375368 359332 375420
rect 359556 375368 359608 375420
rect 218980 372580 219032 372632
rect 219164 372580 219216 372632
rect 218980 367752 219032 367804
rect 219164 367752 219216 367804
rect 359280 365687 359332 365696
rect 359280 365653 359289 365687
rect 359289 365653 359323 365687
rect 359323 365653 359332 365687
rect 359280 365644 359332 365653
rect 364340 364352 364392 364404
rect 364524 364352 364576 364404
rect 218980 360204 219032 360256
rect 359188 360068 359240 360120
rect 218796 354807 218848 354816
rect 218796 354773 218805 354807
rect 218805 354773 218839 354807
rect 218839 354773 218848 354807
rect 218796 354764 218848 354773
rect 218796 354628 218848 354680
rect 218980 350455 219032 350464
rect 218980 350421 218989 350455
rect 218989 350421 219023 350455
rect 219023 350421 219032 350455
rect 218980 350412 219032 350421
rect 364340 345040 364392 345092
rect 364524 345040 364576 345092
rect 218980 340892 219032 340944
rect 218888 340824 218940 340876
rect 3516 338036 3568 338088
rect 352012 338036 352064 338088
rect 3424 337968 3476 338020
rect 270776 337968 270828 338020
rect 286968 337968 287020 338020
rect 363604 337968 363656 338020
rect 238300 337900 238352 337952
rect 359464 337900 359516 337952
rect 254492 337832 254544 337884
rect 364340 337832 364392 337884
rect 218888 337764 218940 337816
rect 303252 337764 303304 337816
rect 319536 337764 319588 337816
rect 366364 337764 366416 337816
rect 3700 337356 3752 337408
rect 335728 337356 335780 337408
rect 358820 335316 358872 335368
rect 359096 335316 359148 335368
rect 358820 325592 358872 325644
rect 359096 325592 359148 325644
rect 358820 316004 358872 316056
rect 359096 316004 359148 316056
rect 358820 306280 358872 306332
rect 359096 306280 359148 306332
rect 358820 296692 358872 296744
rect 359096 296692 359148 296744
rect 358820 286968 358872 287020
rect 359096 286968 359148 287020
rect 3424 280100 3476 280152
rect 358912 280100 358964 280152
rect 358820 277380 358872 277432
rect 359096 277380 359148 277432
rect 358820 267724 358872 267776
rect 359004 267724 359056 267776
rect 358912 260788 358964 260840
rect 358820 251243 358872 251252
rect 358820 251209 358829 251243
rect 358829 251209 358863 251243
rect 358863 251209 358872 251243
rect 358820 251200 358872 251209
rect 358912 241451 358964 241460
rect 358912 241417 358921 241451
rect 358921 241417 358955 241451
rect 358955 241417 358964 241451
rect 358912 241408 358964 241417
rect 359096 234608 359148 234660
rect 358912 222164 358964 222216
rect 359188 222164 359240 222216
rect 359188 215364 359240 215416
rect 359096 215228 359148 215280
rect 358912 202852 358964 202904
rect 359188 202852 359240 202904
rect 359188 196052 359240 196104
rect 359096 195916 359148 195968
rect 358912 183540 358964 183592
rect 359188 183540 359240 183592
rect 359004 173884 359056 173936
rect 359188 173884 359240 173936
rect 358820 151784 358872 151836
rect 359004 151784 359056 151836
rect 358820 132472 358872 132524
rect 359004 132472 359056 132524
rect 358820 113160 358872 113212
rect 359004 113160 359056 113212
rect 358820 93848 358872 93900
rect 359004 93848 359056 93900
rect 358820 74536 358872 74588
rect 359004 74536 359056 74588
rect 358820 55224 358872 55276
rect 359004 55224 359056 55276
rect 358820 35912 358872 35964
rect 359004 35912 359056 35964
rect 358820 16600 358872 16652
rect 359004 16600 359056 16652
rect 572 3408 624 3460
rect 359004 3408 359056 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 154132 695570 154160 703520
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 154224 688634 154252 695506
rect 218992 694210 219020 703520
rect 229008 700528 229060 700534
rect 229008 700470 229060 700476
rect 218980 694204 219032 694210
rect 218980 694146 219032 694152
rect 219164 694204 219216 694210
rect 219164 694146 219216 694152
rect 219176 688702 219204 694146
rect 219164 688696 219216 688702
rect 219164 688638 219216 688644
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 219072 688628 219124 688634
rect 219072 688570 219124 688576
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 219084 678994 219112 688570
rect 218992 678966 219112 678994
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3330 567352 3386 567361
rect 3330 567287 3386 567296
rect 3344 567254 3372 567287
rect 3332 567248 3384 567254
rect 3332 567190 3384 567196
rect 3330 495544 3386 495553
rect 3330 495479 3332 495488
rect 3384 495479 3386 495488
rect 3332 495450 3384 495456
rect 3332 396024 3384 396030
rect 3332 395966 3384 395972
rect 3344 395049 3372 395966
rect 3330 395040 3386 395049
rect 3330 394975 3386 394984
rect 3436 338026 3464 667927
rect 154500 663762 154528 673474
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 154316 663734 154528 663762
rect 154316 654158 154344 663734
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 154500 644450 154528 654094
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 154316 644422 154528 644450
rect 154316 634846 154344 644422
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 154500 625138 154528 634782
rect 219176 630578 219204 637502
rect 219176 630550 219388 630578
rect 219360 626550 219388 630550
rect 219348 626544 219400 626550
rect 219348 626486 219400 626492
rect 154316 625110 154528 625138
rect 3514 624880 3570 624889
rect 3514 624815 3570 624824
rect 3528 338094 3556 624815
rect 154316 615534 154344 625110
rect 219348 616888 219400 616894
rect 219348 616830 219400 616836
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 154500 605826 154528 615470
rect 219360 611454 219388 616830
rect 219348 611448 219400 611454
rect 219348 611390 219400 611396
rect 219072 608728 219124 608734
rect 219072 608670 219124 608676
rect 219084 608598 219112 608670
rect 219072 608592 219124 608598
rect 219072 608534 219124 608540
rect 154316 605798 154528 605826
rect 154316 596222 154344 605798
rect 219256 601588 219308 601594
rect 219256 601530 219308 601536
rect 219268 598942 219296 601530
rect 219256 598936 219308 598942
rect 219256 598878 219308 598884
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 154408 596142 154528 596158
rect 154408 591954 154436 596142
rect 154316 591926 154436 591954
rect 154316 589286 154344 591926
rect 219164 589348 219216 589354
rect 219164 589290 219216 589296
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 219176 582418 219204 589290
rect 218980 582412 219032 582418
rect 218980 582354 219032 582360
rect 219164 582412 219216 582418
rect 219164 582354 219216 582360
rect 154304 579760 154356 579766
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 154224 579686 154344 579702
rect 154224 579630 154252 579686
rect 218992 579630 219020 582354
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 218980 579624 219032 579630
rect 218980 579566 219032 579572
rect 154408 562970 154436 579566
rect 218888 569968 218940 569974
rect 218888 569910 218940 569916
rect 218900 563106 218928 569910
rect 218888 563100 218940 563106
rect 218888 563042 218940 563048
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 218980 562964 219032 562970
rect 218980 562906 219032 562912
rect 154224 553330 154252 562906
rect 218992 560266 219020 562906
rect 218900 560238 219020 560266
rect 218900 553450 218928 560238
rect 218888 553444 218940 553450
rect 218888 553386 218940 553392
rect 154224 553302 154344 553330
rect 154316 543810 154344 553302
rect 218888 550656 218940 550662
rect 218888 550598 218940 550604
rect 154316 543782 154528 543810
rect 218900 543794 218928 550598
rect 154500 534018 154528 543782
rect 218888 543788 218940 543794
rect 218888 543730 218940 543736
rect 218980 543652 219032 543658
rect 218980 543594 219032 543600
rect 218992 540977 219020 543594
rect 218978 540968 219034 540977
rect 218978 540903 219034 540912
rect 219162 540968 219218 540977
rect 219162 540903 219218 540912
rect 154408 533990 154528 534018
rect 154408 531282 154436 533990
rect 219176 533882 219204 540903
rect 218992 533854 219204 533882
rect 218992 531321 219020 533854
rect 218978 531312 219034 531321
rect 154396 531276 154448 531282
rect 218978 531247 219034 531256
rect 219162 531312 219218 531321
rect 219162 531247 219218 531256
rect 154396 531218 154448 531224
rect 219176 524346 219204 531247
rect 218980 524340 219032 524346
rect 218980 524282 219032 524288
rect 219164 524340 219216 524346
rect 219164 524282 219216 524288
rect 154488 521688 154540 521694
rect 154488 521630 154540 521636
rect 154500 514706 154528 521630
rect 154408 514678 154528 514706
rect 218992 514706 219020 524282
rect 218992 514678 219112 514706
rect 154408 511970 154436 514678
rect 219084 512009 219112 514678
rect 218886 512000 218942 512009
rect 154396 511964 154448 511970
rect 218886 511935 218942 511944
rect 219070 512000 219126 512009
rect 219070 511935 219126 511944
rect 154396 511906 154448 511912
rect 218900 502382 218928 511935
rect 154488 502376 154540 502382
rect 154488 502318 154540 502324
rect 218888 502376 218940 502382
rect 218888 502318 218940 502324
rect 219348 502376 219400 502382
rect 219348 502318 219400 502324
rect 154500 495394 154528 502318
rect 219360 495394 219388 502318
rect 154316 495366 154528 495394
rect 219268 495366 219388 495394
rect 154316 485858 154344 495366
rect 219268 485874 219296 495366
rect 154304 485852 154356 485858
rect 154304 485794 154356 485800
rect 219176 485846 219296 485874
rect 154396 485716 154448 485722
rect 154396 485658 154448 485664
rect 154408 483002 154436 485658
rect 154120 482996 154172 483002
rect 154120 482938 154172 482944
rect 154396 482996 154448 483002
rect 154396 482938 154448 482944
rect 154132 473385 154160 482938
rect 219176 480282 219204 485846
rect 219164 480276 219216 480282
rect 219164 480218 219216 480224
rect 219348 480276 219400 480282
rect 219348 480218 219400 480224
rect 219360 480162 219388 480218
rect 219268 480134 219388 480162
rect 154118 473376 154174 473385
rect 154118 473311 154174 473320
rect 154302 473376 154358 473385
rect 154302 473311 154358 473320
rect 154316 472666 154344 473311
rect 154304 472660 154356 472666
rect 154304 472602 154356 472608
rect 3608 472116 3660 472122
rect 3608 472058 3660 472064
rect 3516 338088 3568 338094
rect 3516 338030 3568 338036
rect 3424 338020 3476 338026
rect 3424 337962 3476 337968
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 3422 252512 3478 252521
rect 3422 252447 3478 252456
rect 3436 251297 3464 252447
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3620 208185 3648 472058
rect 3700 472048 3752 472054
rect 3700 471990 3752 471996
rect 3712 438025 3740 471990
rect 219268 470642 219296 480134
rect 219176 470614 219296 470642
rect 219176 460970 219204 470614
rect 219164 460964 219216 460970
rect 219164 460906 219216 460912
rect 219348 460964 219400 460970
rect 219348 460906 219400 460912
rect 219360 460850 219388 460906
rect 219268 460822 219388 460850
rect 219268 444378 219296 460822
rect 228362 448352 228418 448361
rect 228362 448287 228418 448296
rect 219256 444372 219308 444378
rect 219256 444314 219308 444320
rect 219440 444372 219492 444378
rect 219440 444314 219492 444320
rect 3698 438016 3754 438025
rect 3698 437951 3754 437960
rect 219452 434761 219480 444314
rect 219162 434752 219218 434761
rect 219162 434687 219218 434696
rect 219438 434752 219494 434761
rect 219438 434687 219494 434696
rect 219176 427854 219204 434687
rect 218980 427848 219032 427854
rect 218980 427790 219032 427796
rect 219164 427848 219216 427854
rect 219164 427790 219216 427796
rect 218992 425066 219020 427790
rect 218704 425060 218756 425066
rect 218704 425002 218756 425008
rect 218980 425060 219032 425066
rect 218980 425002 219032 425008
rect 218716 415449 218744 425002
rect 218702 415440 218758 415449
rect 218702 415375 218758 415384
rect 218886 415440 218942 415449
rect 218886 415375 218942 415384
rect 218900 408542 218928 415375
rect 218888 408536 218940 408542
rect 218888 408478 218940 408484
rect 218980 408400 219032 408406
rect 218980 408342 219032 408348
rect 218992 405686 219020 408342
rect 218980 405680 219032 405686
rect 218980 405622 219032 405628
rect 218888 396092 218940 396098
rect 218888 396034 218940 396040
rect 218900 395978 218928 396034
rect 228376 396030 228404 448287
rect 229020 404977 229048 700470
rect 283852 700466 283880 703520
rect 295248 700596 295300 700602
rect 295248 700538 295300 700544
rect 283840 700460 283892 700466
rect 283840 700402 283892 700408
rect 240048 700392 240100 700398
rect 240048 700334 240100 700340
rect 240060 470098 240088 700334
rect 276480 472660 276532 472666
rect 276480 472602 276532 472608
rect 257896 472116 257948 472122
rect 257896 472058 257948 472064
rect 239876 470070 240088 470098
rect 239876 469826 239904 470070
rect 257908 469948 257936 472058
rect 276492 469948 276520 472602
rect 295260 469962 295288 700538
rect 300136 700534 300164 703520
rect 348804 700602 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 358912 700460 358964 700466
rect 358912 700402 358964 700408
rect 358820 700324 358872 700330
rect 358820 700266 358872 700272
rect 314568 485852 314620 485858
rect 314568 485794 314620 485800
rect 314580 472734 314608 485794
rect 313648 472728 313700 472734
rect 313648 472670 313700 472676
rect 314568 472728 314620 472734
rect 314568 472670 314620 472676
rect 295090 469934 295288 469962
rect 313660 469948 313688 472670
rect 350816 472048 350868 472054
rect 332230 472016 332286 472025
rect 350816 471990 350868 471996
rect 332230 471951 332286 471960
rect 332244 469948 332272 471951
rect 350828 469948 350856 471990
rect 239430 469798 239904 469826
rect 358832 405634 358860 700266
rect 358924 419370 358952 700402
rect 363604 700324 363656 700330
rect 363604 700266 363656 700272
rect 362224 685908 362276 685914
rect 362224 685850 362276 685856
rect 359004 567248 359056 567254
rect 359004 567190 359056 567196
rect 359016 448746 359044 567190
rect 359096 495508 359148 495514
rect 359096 495450 359148 495456
rect 359108 463162 359136 495450
rect 359554 463176 359610 463185
rect 359108 463134 359554 463162
rect 359554 463111 359610 463120
rect 359554 448760 359610 448769
rect 359016 448718 359554 448746
rect 359554 448695 359610 448704
rect 359464 438932 359516 438938
rect 359464 438874 359516 438880
rect 358924 419354 359228 419370
rect 358924 419348 359240 419354
rect 358924 419342 359188 419348
rect 359188 419290 359240 419296
rect 358832 405618 359228 405634
rect 358832 405612 359240 405618
rect 358832 405606 359188 405612
rect 359188 405554 359240 405560
rect 229006 404968 229062 404977
rect 229006 404903 229062 404912
rect 218808 395950 218928 395978
rect 228364 396024 228416 396030
rect 228364 395966 228416 395972
rect 218808 389042 218836 395950
rect 359188 389496 359240 389502
rect 359016 389444 359188 389450
rect 359016 389438 359240 389444
rect 359016 389422 359228 389438
rect 218808 389014 219020 389042
rect 218992 372638 219020 389014
rect 359016 388498 359044 389422
rect 358924 388470 359044 388498
rect 358924 379386 358952 388470
rect 358924 379358 359044 379386
rect 218980 372632 219032 372638
rect 218980 372574 219032 372580
rect 219164 372632 219216 372638
rect 219164 372574 219216 372580
rect 219176 367810 219204 372574
rect 359016 369866 359044 379358
rect 359280 375420 359332 375426
rect 359280 375362 359332 375368
rect 359016 369838 359136 369866
rect 218980 367804 219032 367810
rect 218980 367746 219032 367752
rect 219164 367804 219216 367810
rect 219164 367746 219216 367752
rect 218992 360262 219020 367746
rect 359108 364392 359136 369838
rect 359292 365702 359320 375362
rect 359280 365696 359332 365702
rect 359280 365638 359332 365644
rect 358924 364364 359136 364392
rect 218980 360256 219032 360262
rect 218980 360198 219032 360204
rect 218796 354816 218848 354822
rect 218796 354758 218848 354764
rect 218808 354686 218836 354758
rect 218796 354680 218848 354686
rect 358924 354634 358952 364364
rect 359188 360120 359240 360126
rect 218796 354622 218848 354628
rect 358832 354606 358952 354634
rect 359108 360068 359188 360074
rect 359108 360062 359240 360068
rect 359108 360046 359228 360062
rect 358832 351778 358860 354606
rect 358740 351750 358860 351778
rect 218980 350464 219032 350470
rect 218980 350406 219032 350412
rect 358740 350418 358768 351750
rect 218992 340950 219020 350406
rect 358740 350390 358952 350418
rect 218980 340944 219032 340950
rect 218980 340886 219032 340892
rect 218888 340876 218940 340882
rect 218888 340818 218940 340824
rect 218900 337822 218928 340818
rect 238312 337958 238340 340068
rect 238300 337952 238352 337958
rect 238300 337894 238352 337900
rect 254504 337890 254532 340068
rect 270788 338026 270816 340068
rect 286980 338026 287008 340068
rect 270776 338020 270828 338026
rect 270776 337962 270828 337968
rect 286968 338020 287020 338026
rect 286968 337962 287020 337968
rect 254492 337884 254544 337890
rect 254492 337826 254544 337832
rect 303264 337822 303292 340068
rect 319548 337822 319576 340068
rect 218888 337816 218940 337822
rect 218888 337758 218940 337764
rect 303252 337816 303304 337822
rect 303252 337758 303304 337764
rect 319536 337816 319588 337822
rect 319536 337758 319588 337764
rect 335740 337414 335768 340068
rect 352024 338094 352052 340068
rect 352012 338088 352064 338094
rect 352012 338030 352064 338036
rect 3700 337408 3752 337414
rect 3700 337350 3752 337356
rect 335728 337408 335780 337414
rect 335728 337350 335780 337356
rect 3712 323105 3740 337350
rect 358820 335368 358872 335374
rect 358820 335310 358872 335316
rect 358832 325650 358860 335310
rect 358820 325644 358872 325650
rect 358820 325586 358872 325592
rect 3698 323096 3754 323105
rect 3698 323031 3754 323040
rect 358820 316056 358872 316062
rect 358820 315998 358872 316004
rect 358832 306338 358860 315998
rect 358820 306332 358872 306338
rect 358820 306274 358872 306280
rect 358820 296744 358872 296750
rect 358820 296686 358872 296692
rect 358832 287026 358860 296686
rect 358820 287020 358872 287026
rect 358820 286962 358872 286968
rect 358924 280158 358952 350390
rect 359108 335374 359136 360046
rect 359476 337958 359504 438874
rect 362236 433945 362264 685850
rect 362316 592068 362368 592074
rect 362316 592010 362368 592016
rect 362222 433936 362278 433945
rect 362222 433871 362278 433880
rect 359556 419348 359608 419354
rect 359556 419290 359608 419296
rect 359568 419257 359596 419290
rect 359554 419248 359610 419257
rect 359554 419183 359610 419192
rect 359556 405612 359608 405618
rect 359556 405554 359608 405560
rect 359568 405521 359596 405554
rect 359554 405512 359610 405521
rect 359554 405447 359610 405456
rect 359554 390008 359610 390017
rect 359554 389943 359610 389952
rect 359568 389502 359596 389943
rect 359556 389496 359608 389502
rect 359556 389438 359608 389444
rect 359554 375592 359610 375601
rect 359554 375527 359610 375536
rect 359568 375426 359596 375527
rect 359556 375420 359608 375426
rect 359556 375362 359608 375368
rect 362328 347313 362356 592010
rect 362408 545148 362460 545154
rect 362408 545090 362460 545096
rect 362420 361729 362448 545090
rect 362406 361720 362462 361729
rect 362406 361655 362462 361664
rect 362314 347304 362370 347313
rect 362314 347239 362370 347248
rect 363616 338026 363644 700266
rect 365088 692850 365116 703446
rect 413664 700466 413692 703520
rect 366364 700460 366416 700466
rect 366364 700402 366416 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 364340 692844 364392 692850
rect 364340 692786 364392 692792
rect 365076 692844 365128 692850
rect 365076 692786 365128 692792
rect 364352 683074 364380 692786
rect 364352 683046 364564 683074
rect 364536 673538 364564 683046
rect 364340 673532 364392 673538
rect 364340 673474 364392 673480
rect 364524 673532 364576 673538
rect 364524 673474 364576 673480
rect 364352 663762 364380 673474
rect 364352 663734 364564 663762
rect 364536 654158 364564 663734
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 364352 644450 364380 654094
rect 364352 644422 364564 644450
rect 364536 634846 364564 644422
rect 364340 634840 364392 634846
rect 364340 634782 364392 634788
rect 364524 634840 364576 634846
rect 364524 634782 364576 634788
rect 364352 625138 364380 634782
rect 364352 625110 364564 625138
rect 364536 615534 364564 625110
rect 364340 615528 364392 615534
rect 364340 615470 364392 615476
rect 364524 615528 364576 615534
rect 364524 615470 364576 615476
rect 364352 605826 364380 615470
rect 364352 605798 364564 605826
rect 364536 596222 364564 605798
rect 364340 596216 364392 596222
rect 364524 596216 364576 596222
rect 364392 596164 364472 596170
rect 364340 596158 364472 596164
rect 364524 596158 364576 596164
rect 364352 596142 364472 596158
rect 364444 596034 364472 596142
rect 364444 596006 364564 596034
rect 364536 591954 364564 596006
rect 364444 591926 364564 591954
rect 364444 589286 364472 591926
rect 364432 589280 364484 589286
rect 364432 589222 364484 589228
rect 364340 579692 364392 579698
rect 364340 579634 364392 579640
rect 364352 572642 364380 579634
rect 364352 572614 364472 572642
rect 364444 569906 364472 572614
rect 364432 569900 364484 569906
rect 364432 569842 364484 569848
rect 364616 563100 364668 563106
rect 364616 563042 364668 563048
rect 364628 560289 364656 563042
rect 364430 560280 364486 560289
rect 364430 560215 364486 560224
rect 364614 560280 364670 560289
rect 364614 560215 364670 560224
rect 364444 550662 364472 560215
rect 364432 550656 364484 550662
rect 364432 550598 364484 550604
rect 364708 550656 364760 550662
rect 364708 550598 364760 550604
rect 364720 543862 364748 550598
rect 364708 543856 364760 543862
rect 364708 543798 364760 543804
rect 364616 543720 364668 543726
rect 364616 543662 364668 543668
rect 364628 540977 364656 543662
rect 364430 540968 364486 540977
rect 364430 540903 364486 540912
rect 364614 540968 364670 540977
rect 364614 540903 364670 540912
rect 364444 531350 364472 540903
rect 364432 531344 364484 531350
rect 364432 531286 364484 531292
rect 364708 531344 364760 531350
rect 364708 531286 364760 531292
rect 364720 524550 364748 531286
rect 364708 524544 364760 524550
rect 364708 524486 364760 524492
rect 364616 524408 364668 524414
rect 364616 524350 364668 524356
rect 364628 521665 364656 524350
rect 364430 521656 364486 521665
rect 364430 521591 364486 521600
rect 364614 521656 364670 521665
rect 364614 521591 364670 521600
rect 364444 512038 364472 521591
rect 364432 512032 364484 512038
rect 364432 511974 364484 511980
rect 364708 512032 364760 512038
rect 364708 511974 364760 511980
rect 364720 502382 364748 511974
rect 364524 502376 364576 502382
rect 364246 502344 364302 502353
rect 364246 502279 364302 502288
rect 364522 502344 364524 502353
rect 364708 502376 364760 502382
rect 364576 502344 364578 502353
rect 364708 502318 364760 502324
rect 364522 502279 364578 502288
rect 364260 492697 364288 502279
rect 364246 492688 364302 492697
rect 364246 492623 364302 492632
rect 364430 492688 364486 492697
rect 364430 492623 364486 492632
rect 364444 489954 364472 492623
rect 364444 489926 364564 489954
rect 364536 480282 364564 489926
rect 364340 480276 364392 480282
rect 364340 480218 364392 480224
rect 364524 480276 364576 480282
rect 364524 480218 364576 480224
rect 364352 480162 364380 480218
rect 364352 480134 364472 480162
rect 364444 470642 364472 480134
rect 364444 470614 364564 470642
rect 364536 460970 364564 470614
rect 364340 460964 364392 460970
rect 364340 460906 364392 460912
rect 364524 460964 364576 460970
rect 364524 460906 364576 460912
rect 364352 460850 364380 460906
rect 364352 460822 364472 460850
rect 364444 451330 364472 460822
rect 364444 451302 364564 451330
rect 364536 441658 364564 451302
rect 364340 441652 364392 441658
rect 364340 441594 364392 441600
rect 364524 441652 364576 441658
rect 364524 441594 364576 441600
rect 364352 441538 364380 441594
rect 364352 441510 364472 441538
rect 364444 432018 364472 441510
rect 364444 431990 364564 432018
rect 364536 422346 364564 431990
rect 364340 422340 364392 422346
rect 364340 422282 364392 422288
rect 364524 422340 364576 422346
rect 364524 422282 364576 422288
rect 364352 422226 364380 422282
rect 364352 422198 364472 422226
rect 364444 412706 364472 422198
rect 364444 412678 364564 412706
rect 364536 403034 364564 412678
rect 364340 403028 364392 403034
rect 364340 402970 364392 402976
rect 364524 403028 364576 403034
rect 364524 402970 364576 402976
rect 364352 402914 364380 402970
rect 364352 402886 364472 402914
rect 364444 393394 364472 402886
rect 364444 393366 364564 393394
rect 364536 383722 364564 393366
rect 364340 383716 364392 383722
rect 364340 383658 364392 383664
rect 364524 383716 364576 383722
rect 364524 383658 364576 383664
rect 364352 383602 364380 383658
rect 364352 383574 364472 383602
rect 364444 374082 364472 383574
rect 364444 374054 364564 374082
rect 364536 364410 364564 374054
rect 364340 364404 364392 364410
rect 364340 364346 364392 364352
rect 364524 364404 364576 364410
rect 364524 364346 364576 364352
rect 364352 354634 364380 364346
rect 364352 354606 364564 354634
rect 364536 345098 364564 354606
rect 364340 345092 364392 345098
rect 364340 345034 364392 345040
rect 364524 345092 364576 345098
rect 364524 345034 364576 345040
rect 363604 338020 363656 338026
rect 363604 337962 363656 337968
rect 359464 337952 359516 337958
rect 359464 337894 359516 337900
rect 364352 337890 364380 345034
rect 364340 337884 364392 337890
rect 364340 337826 364392 337832
rect 366376 337822 366404 700402
rect 478524 700330 478552 703520
rect 543476 700398 543504 703520
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 478512 700324 478564 700330
rect 478512 700266 478564 700272
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 580262 393000 580318 393009
rect 580262 392935 580318 392944
rect 580276 362953 580304 392935
rect 580262 362944 580318 362953
rect 580262 362879 580318 362888
rect 366364 337816 366416 337822
rect 366364 337758 366416 337764
rect 359096 335368 359148 335374
rect 359096 335310 359148 335316
rect 359096 325644 359148 325650
rect 359096 325586 359148 325592
rect 359108 316062 359136 325586
rect 359096 316056 359148 316062
rect 359096 315998 359148 316004
rect 359096 306332 359148 306338
rect 359096 306274 359148 306280
rect 359108 296750 359136 306274
rect 359096 296744 359148 296750
rect 359096 296686 359148 296692
rect 359096 287020 359148 287026
rect 359096 286962 359148 286968
rect 358912 280152 358964 280158
rect 358912 280094 358964 280100
rect 358832 277438 358860 277469
rect 359108 277438 359136 286962
rect 358820 277432 358872 277438
rect 359096 277432 359148 277438
rect 358872 277380 359044 277386
rect 358820 277374 359044 277380
rect 359096 277374 359148 277380
rect 358832 277358 359044 277374
rect 359016 267782 359044 277358
rect 358820 267776 358872 267782
rect 359004 267776 359056 267782
rect 358872 267724 358952 267730
rect 358820 267718 358952 267724
rect 359004 267718 359056 267724
rect 358832 267702 358952 267718
rect 358924 267594 358952 267702
rect 358924 267566 359044 267594
rect 359016 263514 359044 267566
rect 358924 263486 359044 263514
rect 358924 260846 358952 263486
rect 358912 260840 358964 260846
rect 358912 260782 358964 260788
rect 358820 251252 358872 251258
rect 358820 251194 358872 251200
rect 358832 244202 358860 251194
rect 358832 244174 358952 244202
rect 358924 241466 358952 244174
rect 358912 241460 358964 241466
rect 358912 241402 358964 241408
rect 359096 234660 359148 234666
rect 359096 234602 359148 234608
rect 359108 231849 359136 234602
rect 358910 231840 358966 231849
rect 358910 231775 358966 231784
rect 359094 231840 359150 231849
rect 359094 231775 359150 231784
rect 358924 222222 358952 231775
rect 358912 222216 358964 222222
rect 358912 222158 358964 222164
rect 359188 222216 359240 222222
rect 359188 222158 359240 222164
rect 359200 215422 359228 222158
rect 359188 215416 359240 215422
rect 359188 215358 359240 215364
rect 359096 215280 359148 215286
rect 359096 215222 359148 215228
rect 359108 212537 359136 215222
rect 358910 212528 358966 212537
rect 358910 212463 358966 212472
rect 359094 212528 359150 212537
rect 359094 212463 359150 212472
rect 3606 208176 3662 208185
rect 3606 208111 3662 208120
rect 358924 202910 358952 212463
rect 358912 202904 358964 202910
rect 358912 202846 358964 202852
rect 359188 202904 359240 202910
rect 359188 202846 359240 202852
rect 359200 196110 359228 202846
rect 359188 196104 359240 196110
rect 359188 196046 359240 196052
rect 359096 195968 359148 195974
rect 359096 195910 359148 195916
rect 359108 193225 359136 195910
rect 358910 193216 358966 193225
rect 358910 193151 358966 193160
rect 359094 193216 359150 193225
rect 359094 193151 359150 193160
rect 358924 183598 358952 193151
rect 358912 183592 358964 183598
rect 358912 183534 358964 183540
rect 359188 183592 359240 183598
rect 359188 183534 359240 183540
rect 359200 173942 359228 183534
rect 359004 173936 359056 173942
rect 358726 173904 358782 173913
rect 358726 173839 358782 173848
rect 359002 173904 359004 173913
rect 359188 173936 359240 173942
rect 359056 173904 359058 173913
rect 359188 173878 359240 173884
rect 359002 173839 359058 173848
rect 358740 164257 358768 173839
rect 358726 164248 358782 164257
rect 358726 164183 358782 164192
rect 358910 164248 358966 164257
rect 358910 164183 358966 164192
rect 358924 161514 358952 164183
rect 358924 161486 359044 161514
rect 359016 151842 359044 161486
rect 358820 151836 358872 151842
rect 358820 151778 358872 151784
rect 359004 151836 359056 151842
rect 359004 151778 359056 151784
rect 358832 151722 358860 151778
rect 358832 151694 358952 151722
rect 358924 142202 358952 151694
rect 358924 142174 359044 142202
rect 359016 132530 359044 142174
rect 358820 132524 358872 132530
rect 358820 132466 358872 132472
rect 359004 132524 359056 132530
rect 359004 132466 359056 132472
rect 358832 132410 358860 132466
rect 358832 132382 358952 132410
rect 358924 122890 358952 132382
rect 358924 122862 359044 122890
rect 359016 113218 359044 122862
rect 358820 113212 358872 113218
rect 358820 113154 358872 113160
rect 359004 113212 359056 113218
rect 359004 113154 359056 113160
rect 358832 113098 358860 113154
rect 358832 113070 358952 113098
rect 358924 103578 358952 113070
rect 358924 103550 359044 103578
rect 359016 93906 359044 103550
rect 358820 93900 358872 93906
rect 358820 93842 358872 93848
rect 359004 93900 359056 93906
rect 359004 93842 359056 93848
rect 358832 93786 358860 93842
rect 358832 93758 358952 93786
rect 358924 84266 358952 93758
rect 358924 84238 359044 84266
rect 359016 74594 359044 84238
rect 358820 74588 358872 74594
rect 358820 74530 358872 74536
rect 359004 74588 359056 74594
rect 359004 74530 359056 74536
rect 358832 74474 358860 74530
rect 358832 74446 358952 74474
rect 358924 64954 358952 74446
rect 358924 64926 359044 64954
rect 359016 55282 359044 64926
rect 358820 55276 358872 55282
rect 358820 55218 358872 55224
rect 359004 55276 359056 55282
rect 359004 55218 359056 55224
rect 358832 55162 358860 55218
rect 358832 55134 358952 55162
rect 358924 45642 358952 55134
rect 358924 45614 359044 45642
rect 359016 35970 359044 45614
rect 358820 35964 358872 35970
rect 358820 35906 358872 35912
rect 359004 35964 359056 35970
rect 359004 35906 359056 35912
rect 358832 26194 358860 35906
rect 358832 26166 359044 26194
rect 359016 16658 359044 26166
rect 358820 16652 358872 16658
rect 358820 16594 358872 16600
rect 359004 16652 359056 16658
rect 359004 16594 359056 16600
rect 358832 6882 358860 16594
rect 358832 6854 359044 6882
rect 359016 3466 359044 6854
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 359004 3460 359056 3466
rect 359004 3402 359056 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 667936 3478 667992
rect 3330 567296 3386 567352
rect 3330 495508 3386 495544
rect 3330 495488 3332 495508
rect 3332 495488 3384 495508
rect 3384 495488 3386 495508
rect 3330 394984 3386 395040
rect 3514 624824 3570 624880
rect 218978 540912 219034 540968
rect 219162 540912 219218 540968
rect 218978 531256 219034 531312
rect 219162 531256 219218 531312
rect 218886 511944 218942 512000
rect 219070 511944 219126 512000
rect 154118 473320 154174 473376
rect 154302 473320 154358 473376
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 3422 252456 3478 252512
rect 3422 251232 3478 251288
rect 228362 448296 228418 448352
rect 3698 437960 3754 438016
rect 219162 434696 219218 434752
rect 219438 434696 219494 434752
rect 218702 415384 218758 415440
rect 218886 415384 218942 415440
rect 332230 471960 332286 472016
rect 359554 463120 359610 463176
rect 359554 448704 359610 448760
rect 229006 404912 229062 404968
rect 3698 323040 3754 323096
rect 362222 433880 362278 433936
rect 359554 419192 359610 419248
rect 359554 405456 359610 405512
rect 359554 389952 359610 390008
rect 359554 375536 359610 375592
rect 362406 361664 362462 361720
rect 362314 347248 362370 347304
rect 364430 560224 364486 560280
rect 364614 560224 364670 560280
rect 364430 540912 364486 540968
rect 364614 540912 364670 540968
rect 364430 521600 364486 521656
rect 364614 521600 364670 521656
rect 364246 502288 364302 502344
rect 364522 502324 364524 502344
rect 364524 502324 364576 502344
rect 364576 502324 364578 502344
rect 364522 502288 364578 502324
rect 364246 492632 364302 492688
rect 364430 492632 364486 492688
rect 580170 686296 580226 686352
rect 580170 592456 580226 592512
rect 580170 545536 580226 545592
rect 580170 486784 580226 486840
rect 580170 439864 580226 439920
rect 580262 392944 580318 393000
rect 580262 362888 580318 362944
rect 358910 231784 358966 231840
rect 359094 231784 359150 231840
rect 358910 212472 358966 212528
rect 359094 212472 359150 212528
rect 3606 208120 3662 208176
rect 358910 193160 358966 193216
rect 359094 193160 359150 193216
rect 358726 173848 358782 173904
rect 359002 173884 359004 173904
rect 359004 173884 359056 173904
rect 359056 173884 359058 173904
rect 359002 173848 359058 173884
rect 358726 164192 358782 164248
rect 358910 164192 358966 164248
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653428 480 653668
rect 583520 650980 584960 651220
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 583520 627588 584960 627828
rect -960 624882 480 624972
rect 3509 624882 3575 624885
rect -960 624880 3575 624882
rect -960 624824 3514 624880
rect 3570 624824 3575 624880
rect -960 624822 3575 624824
rect -960 624732 480 624822
rect 3509 624819 3575 624822
rect 583520 615756 584960 615996
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 583520 580668 584960 580908
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3325 567354 3391 567357
rect -960 567352 3391 567354
rect -960 567296 3330 567352
rect 3386 567296 3391 567352
rect -960 567294 3391 567296
rect -960 567204 480 567294
rect 3325 567291 3391 567294
rect 364425 560282 364491 560285
rect 364609 560282 364675 560285
rect 364425 560280 364675 560282
rect 364425 560224 364430 560280
rect 364486 560224 364614 560280
rect 364670 560224 364675 560280
rect 364425 560222 364675 560224
rect 364425 560219 364491 560222
rect 364609 560219 364675 560222
rect 583520 557140 584960 557380
rect -960 552924 480 553164
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 218973 540970 219039 540973
rect 219157 540970 219223 540973
rect 218973 540968 219223 540970
rect 218973 540912 218978 540968
rect 219034 540912 219162 540968
rect 219218 540912 219223 540968
rect 218973 540910 219223 540912
rect 218973 540907 219039 540910
rect 219157 540907 219223 540910
rect 364425 540970 364491 540973
rect 364609 540970 364675 540973
rect 364425 540968 364675 540970
rect 364425 540912 364430 540968
rect 364486 540912 364614 540968
rect 364670 540912 364675 540968
rect 364425 540910 364675 540912
rect 364425 540907 364491 540910
rect 364609 540907 364675 540910
rect -960 538508 480 538748
rect 583520 533748 584960 533988
rect 218973 531314 219039 531317
rect 219157 531314 219223 531317
rect 218973 531312 219223 531314
rect 218973 531256 218978 531312
rect 219034 531256 219162 531312
rect 219218 531256 219223 531312
rect 218973 531254 219223 531256
rect 218973 531251 219039 531254
rect 219157 531251 219223 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 364425 521658 364491 521661
rect 364609 521658 364675 521661
rect 364425 521656 364675 521658
rect 364425 521600 364430 521656
rect 364486 521600 364614 521656
rect 364670 521600 364675 521656
rect 364425 521598 364675 521600
rect 364425 521595 364491 521598
rect 364609 521595 364675 521598
rect 218881 512002 218947 512005
rect 219065 512002 219131 512005
rect 218881 512000 219131 512002
rect 218881 511944 218886 512000
rect 218942 511944 219070 512000
rect 219126 511944 219131 512000
rect 218881 511942 219131 511944
rect 218881 511939 218947 511942
rect 219065 511939 219131 511942
rect 583520 510220 584960 510460
rect -960 509812 480 510052
rect 364241 502346 364307 502349
rect 364517 502346 364583 502349
rect 364241 502344 364583 502346
rect 364241 502288 364246 502344
rect 364302 502288 364522 502344
rect 364578 502288 364583 502344
rect 364241 502286 364583 502288
rect 364241 502283 364307 502286
rect 364517 502283 364583 502286
rect 583520 498524 584960 498764
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 364241 492690 364307 492693
rect 364425 492690 364491 492693
rect 364241 492688 364491 492690
rect 364241 492632 364246 492688
rect 364302 492632 364430 492688
rect 364486 492632 364491 492688
rect 364241 492630 364491 492632
rect 364241 492627 364307 492630
rect 364425 492627 364491 492630
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect -960 480980 480 481220
rect 583520 474996 584960 475236
rect 154113 473378 154179 473381
rect 154297 473378 154363 473381
rect 154113 473376 154363 473378
rect 154113 473320 154118 473376
rect 154174 473320 154302 473376
rect 154358 473320 154363 473376
rect 154113 473318 154363 473320
rect 154113 473315 154179 473318
rect 154297 473315 154363 473318
rect 268326 471956 268332 472020
rect 268396 472018 268402 472020
rect 332225 472018 332291 472021
rect 268396 472016 332291 472018
rect 268396 471960 332230 472016
rect 332286 471960 332291 472016
rect 268396 471958 332291 471960
rect 268396 471956 268402 471958
rect 332225 471955 332291 471958
rect -960 466700 480 466940
rect 583520 463300 584960 463540
rect 359549 463178 359615 463181
rect 359549 463176 359658 463178
rect 359549 463120 359554 463176
rect 359610 463120 359658 463176
rect 359549 463115 359658 463120
rect 359598 462740 359658 463115
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 359549 448762 359615 448765
rect 359549 448760 359658 448762
rect 359549 448704 359554 448760
rect 359610 448704 359658 448760
rect 359549 448699 359658 448704
rect 228357 448354 228423 448357
rect 228357 448352 230276 448354
rect 228357 448296 228362 448352
rect 228418 448296 230276 448352
rect 359598 448324 359658 448699
rect 228357 448294 230276 448296
rect 228357 448291 228423 448294
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3693 438018 3759 438021
rect -960 438016 3759 438018
rect -960 437960 3698 438016
rect 3754 437960 3759 438016
rect -960 437958 3759 437960
rect -960 437868 480 437958
rect 3693 437955 3759 437958
rect 219157 434754 219223 434757
rect 219433 434754 219499 434757
rect 219157 434752 219499 434754
rect 219157 434696 219162 434752
rect 219218 434696 219438 434752
rect 219494 434696 219499 434752
rect 219157 434694 219499 434696
rect 219157 434691 219223 434694
rect 219433 434691 219499 434694
rect 362217 433938 362283 433941
rect 360180 433936 362283 433938
rect 360180 433880 362222 433936
rect 362278 433880 362283 433936
rect 360180 433878 362283 433880
rect 362217 433875 362283 433878
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 359598 419253 359658 419492
rect 359549 419248 359658 419253
rect 359549 419192 359554 419248
rect 359610 419192 359658 419248
rect 359549 419190 359658 419192
rect 359549 419187 359615 419190
rect 583520 416380 584960 416620
rect 218697 415442 218763 415445
rect 218881 415442 218947 415445
rect 218697 415440 218947 415442
rect 218697 415384 218702 415440
rect 218758 415384 218886 415440
rect 218942 415384 218947 415440
rect 218697 415382 218947 415384
rect 218697 415379 218763 415382
rect 218881 415379 218947 415382
rect -960 409172 480 409412
rect 359549 405514 359615 405517
rect 359549 405512 359658 405514
rect 359549 405456 359554 405512
rect 359610 405456 359658 405512
rect 359549 405451 359658 405456
rect 229001 404970 229067 404973
rect 229001 404968 230276 404970
rect 229001 404912 229006 404968
rect 229062 404912 230276 404968
rect 359598 404940 359658 405451
rect 229001 404910 230276 404912
rect 229001 404907 229067 404910
rect 583520 404684 584960 404924
rect -960 395042 480 395132
rect 3325 395042 3391 395045
rect -960 395040 3391 395042
rect -960 394984 3330 395040
rect 3386 394984 3391 395040
rect -960 394982 3391 394984
rect -960 394892 480 394982
rect 3325 394979 3391 394982
rect 580257 393002 580323 393005
rect 583520 393002 584960 393092
rect 580257 393000 584960 393002
rect 580257 392944 580262 393000
rect 580318 392944 584960 393000
rect 580257 392942 584960 392944
rect 580257 392939 580323 392942
rect 583520 392852 584960 392942
rect 359598 390013 359658 390524
rect 359549 390008 359658 390013
rect 359549 389952 359554 390008
rect 359610 389952 359658 390008
rect 359549 389950 359658 389952
rect 359549 389947 359615 389950
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 359598 375597 359658 376108
rect 359549 375592 359658 375597
rect 359549 375536 359554 375592
rect 359610 375536 359658 375592
rect 359549 375534 359658 375536
rect 359549 375531 359615 375534
rect 583520 369460 584960 369700
rect -960 366060 480 366300
rect 359590 362884 359596 362948
rect 359660 362946 359666 362948
rect 580257 362946 580323 362949
rect 359660 362944 580323 362946
rect 359660 362888 580262 362944
rect 580318 362888 580323 362944
rect 359660 362886 580323 362888
rect 359660 362884 359666 362886
rect 580257 362883 580323 362886
rect 362401 361722 362467 361725
rect 360180 361720 362467 361722
rect 230798 361180 230858 361692
rect 360180 361664 362406 361720
rect 362462 361664 362467 361720
rect 360180 361662 362467 361664
rect 362401 361659 362467 361662
rect 230790 361116 230796 361180
rect 230860 361116 230866 361180
rect 583520 357764 584960 358004
rect -960 351780 480 352020
rect 362309 347306 362375 347309
rect 360180 347304 362375 347306
rect 360180 347248 362314 347304
rect 362370 347248 362375 347304
rect 360180 347246 362375 347248
rect 362309 347243 362375 347246
rect 583520 345932 584960 346172
rect -960 337364 480 337604
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 3693 323098 3759 323101
rect -960 323096 3759 323098
rect -960 323040 3698 323096
rect 3754 323040 3759 323096
rect -960 323038 3759 323040
rect -960 322948 480 323038
rect 3693 323035 3759 323038
rect 583520 322540 584960 322780
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 583520 275620 584960 275860
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 3417 252514 3483 252517
rect 268326 252514 268332 252516
rect 3417 252512 268332 252514
rect 3417 252456 3422 252512
rect 3478 252456 268332 252512
rect 3417 252454 268332 252456
rect 3417 252451 3483 252454
rect 268326 252452 268332 252454
rect 268396 252452 268402 252516
rect 583520 252092 584960 252332
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 583520 240396 584960 240636
rect -960 236860 480 237100
rect 358905 231842 358971 231845
rect 359089 231842 359155 231845
rect 358905 231840 359155 231842
rect 358905 231784 358910 231840
rect 358966 231784 359094 231840
rect 359150 231784 359155 231840
rect 358905 231782 359155 231784
rect 358905 231779 358971 231782
rect 359089 231779 359155 231782
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect 358905 212530 358971 212533
rect 359089 212530 359155 212533
rect 358905 212528 359155 212530
rect 358905 212472 358910 212528
rect 358966 212472 359094 212528
rect 359150 212472 359155 212528
rect 358905 212470 359155 212472
rect 358905 212467 358971 212470
rect 359089 212467 359155 212470
rect -960 208178 480 208268
rect 3601 208178 3667 208181
rect -960 208176 3667 208178
rect -960 208120 3606 208176
rect 3662 208120 3667 208176
rect -960 208118 3667 208120
rect -960 208028 480 208118
rect 3601 208115 3667 208118
rect 583520 205172 584960 205412
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 358905 193218 358971 193221
rect 359089 193218 359155 193221
rect 358905 193216 359155 193218
rect 358905 193160 358910 193216
rect 358966 193160 359094 193216
rect 359150 193160 359155 193216
rect 358905 193158 359155 193160
rect 358905 193155 358971 193158
rect 359089 193155 359155 193158
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 358721 173906 358787 173909
rect 358997 173906 359063 173909
rect 358721 173904 359063 173906
rect 358721 173848 358726 173904
rect 358782 173848 359002 173904
rect 359058 173848 359063 173904
rect 358721 173846 359063 173848
rect 358721 173843 358787 173846
rect 358997 173843 359063 173846
rect 583520 169948 584960 170188
rect -960 164916 480 165156
rect 358721 164250 358787 164253
rect 358905 164250 358971 164253
rect 358721 164248 358971 164250
rect 358721 164192 358726 164248
rect 358782 164192 358910 164248
rect 358966 164192 358971 164248
rect 358721 164190 358971 164192
rect 358721 164187 358787 164190
rect 358905 164187 358971 164190
rect 583520 158252 584960 158492
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 583520 99636 584960 99876
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 583520 17492 584960 17732
rect -960 7020 480 7260
rect 583520 5796 584960 6036
<< via3 >>
rect 268332 471956 268396 472020
rect 359596 362884 359660 362948
rect 230796 361116 230860 361180
rect 268332 252452 268396 252516
<< metal4 >>
rect -8426 711278 -7846 711290
rect -8426 711042 -8254 711278
rect -8018 711042 -7846 711278
rect -8426 710958 -7846 711042
rect -8426 710722 -8254 710958
rect -8018 710722 -7846 710958
rect -8426 678894 -7846 710722
rect -8426 678658 -8254 678894
rect -8018 678658 -7846 678894
rect -8426 678574 -7846 678658
rect -8426 678338 -8254 678574
rect -8018 678338 -7846 678574
rect -8426 642894 -7846 678338
rect -8426 642658 -8254 642894
rect -8018 642658 -7846 642894
rect -8426 642574 -7846 642658
rect -8426 642338 -8254 642574
rect -8018 642338 -7846 642574
rect -8426 606894 -7846 642338
rect -8426 606658 -8254 606894
rect -8018 606658 -7846 606894
rect -8426 606574 -7846 606658
rect -8426 606338 -8254 606574
rect -8018 606338 -7846 606574
rect -8426 570894 -7846 606338
rect -8426 570658 -8254 570894
rect -8018 570658 -7846 570894
rect -8426 570574 -7846 570658
rect -8426 570338 -8254 570574
rect -8018 570338 -7846 570574
rect -8426 534894 -7846 570338
rect -8426 534658 -8254 534894
rect -8018 534658 -7846 534894
rect -8426 534574 -7846 534658
rect -8426 534338 -8254 534574
rect -8018 534338 -7846 534574
rect -8426 498894 -7846 534338
rect -8426 498658 -8254 498894
rect -8018 498658 -7846 498894
rect -8426 498574 -7846 498658
rect -8426 498338 -8254 498574
rect -8018 498338 -7846 498574
rect -8426 462894 -7846 498338
rect -8426 462658 -8254 462894
rect -8018 462658 -7846 462894
rect -8426 462574 -7846 462658
rect -8426 462338 -8254 462574
rect -8018 462338 -7846 462574
rect -8426 426894 -7846 462338
rect -8426 426658 -8254 426894
rect -8018 426658 -7846 426894
rect -8426 426574 -7846 426658
rect -8426 426338 -8254 426574
rect -8018 426338 -7846 426574
rect -8426 390894 -7846 426338
rect -8426 390658 -8254 390894
rect -8018 390658 -7846 390894
rect -8426 390574 -7846 390658
rect -8426 390338 -8254 390574
rect -8018 390338 -7846 390574
rect -8426 354894 -7846 390338
rect -8426 354658 -8254 354894
rect -8018 354658 -7846 354894
rect -8426 354574 -7846 354658
rect -8426 354338 -8254 354574
rect -8018 354338 -7846 354574
rect -8426 318894 -7846 354338
rect -8426 318658 -8254 318894
rect -8018 318658 -7846 318894
rect -8426 318574 -7846 318658
rect -8426 318338 -8254 318574
rect -8018 318338 -7846 318574
rect -8426 282894 -7846 318338
rect -8426 282658 -8254 282894
rect -8018 282658 -7846 282894
rect -8426 282574 -7846 282658
rect -8426 282338 -8254 282574
rect -8018 282338 -7846 282574
rect -8426 246894 -7846 282338
rect -8426 246658 -8254 246894
rect -8018 246658 -7846 246894
rect -8426 246574 -7846 246658
rect -8426 246338 -8254 246574
rect -8018 246338 -7846 246574
rect -8426 210894 -7846 246338
rect -8426 210658 -8254 210894
rect -8018 210658 -7846 210894
rect -8426 210574 -7846 210658
rect -8426 210338 -8254 210574
rect -8018 210338 -7846 210574
rect -8426 174894 -7846 210338
rect -8426 174658 -8254 174894
rect -8018 174658 -7846 174894
rect -8426 174574 -7846 174658
rect -8426 174338 -8254 174574
rect -8018 174338 -7846 174574
rect -8426 138894 -7846 174338
rect -8426 138658 -8254 138894
rect -8018 138658 -7846 138894
rect -8426 138574 -7846 138658
rect -8426 138338 -8254 138574
rect -8018 138338 -7846 138574
rect -8426 102894 -7846 138338
rect -8426 102658 -8254 102894
rect -8018 102658 -7846 102894
rect -8426 102574 -7846 102658
rect -8426 102338 -8254 102574
rect -8018 102338 -7846 102574
rect -8426 66894 -7846 102338
rect -8426 66658 -8254 66894
rect -8018 66658 -7846 66894
rect -8426 66574 -7846 66658
rect -8426 66338 -8254 66574
rect -8018 66338 -7846 66574
rect -8426 30894 -7846 66338
rect -8426 30658 -8254 30894
rect -8018 30658 -7846 30894
rect -8426 30574 -7846 30658
rect -8426 30338 -8254 30574
rect -8018 30338 -7846 30574
rect -8426 -6786 -7846 30338
rect -7506 710358 -6926 710370
rect -7506 710122 -7334 710358
rect -7098 710122 -6926 710358
rect -7506 710038 -6926 710122
rect -7506 709802 -7334 710038
rect -7098 709802 -6926 710038
rect -7506 696894 -6926 709802
rect 11254 710358 11834 711290
rect 11254 710122 11426 710358
rect 11662 710122 11834 710358
rect 11254 710038 11834 710122
rect 11254 709802 11426 710038
rect 11662 709802 11834 710038
rect -7506 696658 -7334 696894
rect -7098 696658 -6926 696894
rect -7506 696574 -6926 696658
rect -7506 696338 -7334 696574
rect -7098 696338 -6926 696574
rect -7506 660894 -6926 696338
rect -7506 660658 -7334 660894
rect -7098 660658 -6926 660894
rect -7506 660574 -6926 660658
rect -7506 660338 -7334 660574
rect -7098 660338 -6926 660574
rect -7506 624894 -6926 660338
rect -7506 624658 -7334 624894
rect -7098 624658 -6926 624894
rect -7506 624574 -6926 624658
rect -7506 624338 -7334 624574
rect -7098 624338 -6926 624574
rect -7506 588894 -6926 624338
rect -7506 588658 -7334 588894
rect -7098 588658 -6926 588894
rect -7506 588574 -6926 588658
rect -7506 588338 -7334 588574
rect -7098 588338 -6926 588574
rect -7506 552894 -6926 588338
rect -7506 552658 -7334 552894
rect -7098 552658 -6926 552894
rect -7506 552574 -6926 552658
rect -7506 552338 -7334 552574
rect -7098 552338 -6926 552574
rect -7506 516894 -6926 552338
rect -7506 516658 -7334 516894
rect -7098 516658 -6926 516894
rect -7506 516574 -6926 516658
rect -7506 516338 -7334 516574
rect -7098 516338 -6926 516574
rect -7506 480894 -6926 516338
rect -7506 480658 -7334 480894
rect -7098 480658 -6926 480894
rect -7506 480574 -6926 480658
rect -7506 480338 -7334 480574
rect -7098 480338 -6926 480574
rect -7506 444894 -6926 480338
rect -7506 444658 -7334 444894
rect -7098 444658 -6926 444894
rect -7506 444574 -6926 444658
rect -7506 444338 -7334 444574
rect -7098 444338 -6926 444574
rect -7506 408894 -6926 444338
rect -7506 408658 -7334 408894
rect -7098 408658 -6926 408894
rect -7506 408574 -6926 408658
rect -7506 408338 -7334 408574
rect -7098 408338 -6926 408574
rect -7506 372894 -6926 408338
rect -7506 372658 -7334 372894
rect -7098 372658 -6926 372894
rect -7506 372574 -6926 372658
rect -7506 372338 -7334 372574
rect -7098 372338 -6926 372574
rect -7506 336894 -6926 372338
rect -7506 336658 -7334 336894
rect -7098 336658 -6926 336894
rect -7506 336574 -6926 336658
rect -7506 336338 -7334 336574
rect -7098 336338 -6926 336574
rect -7506 300894 -6926 336338
rect -7506 300658 -7334 300894
rect -7098 300658 -6926 300894
rect -7506 300574 -6926 300658
rect -7506 300338 -7334 300574
rect -7098 300338 -6926 300574
rect -7506 264894 -6926 300338
rect -7506 264658 -7334 264894
rect -7098 264658 -6926 264894
rect -7506 264574 -6926 264658
rect -7506 264338 -7334 264574
rect -7098 264338 -6926 264574
rect -7506 228894 -6926 264338
rect -7506 228658 -7334 228894
rect -7098 228658 -6926 228894
rect -7506 228574 -6926 228658
rect -7506 228338 -7334 228574
rect -7098 228338 -6926 228574
rect -7506 192894 -6926 228338
rect -7506 192658 -7334 192894
rect -7098 192658 -6926 192894
rect -7506 192574 -6926 192658
rect -7506 192338 -7334 192574
rect -7098 192338 -6926 192574
rect -7506 156894 -6926 192338
rect -7506 156658 -7334 156894
rect -7098 156658 -6926 156894
rect -7506 156574 -6926 156658
rect -7506 156338 -7334 156574
rect -7098 156338 -6926 156574
rect -7506 120894 -6926 156338
rect -7506 120658 -7334 120894
rect -7098 120658 -6926 120894
rect -7506 120574 -6926 120658
rect -7506 120338 -7334 120574
rect -7098 120338 -6926 120574
rect -7506 84894 -6926 120338
rect -7506 84658 -7334 84894
rect -7098 84658 -6926 84894
rect -7506 84574 -6926 84658
rect -7506 84338 -7334 84574
rect -7098 84338 -6926 84574
rect -7506 48894 -6926 84338
rect -7506 48658 -7334 48894
rect -7098 48658 -6926 48894
rect -7506 48574 -6926 48658
rect -7506 48338 -7334 48574
rect -7098 48338 -6926 48574
rect -7506 12894 -6926 48338
rect -7506 12658 -7334 12894
rect -7098 12658 -6926 12894
rect -7506 12574 -6926 12658
rect -7506 12338 -7334 12574
rect -7098 12338 -6926 12574
rect -7506 -5866 -6926 12338
rect -6586 709438 -6006 709450
rect -6586 709202 -6414 709438
rect -6178 709202 -6006 709438
rect -6586 709118 -6006 709202
rect -6586 708882 -6414 709118
rect -6178 708882 -6006 709118
rect -6586 675414 -6006 708882
rect -6586 675178 -6414 675414
rect -6178 675178 -6006 675414
rect -6586 675094 -6006 675178
rect -6586 674858 -6414 675094
rect -6178 674858 -6006 675094
rect -6586 639414 -6006 674858
rect -6586 639178 -6414 639414
rect -6178 639178 -6006 639414
rect -6586 639094 -6006 639178
rect -6586 638858 -6414 639094
rect -6178 638858 -6006 639094
rect -6586 603414 -6006 638858
rect -6586 603178 -6414 603414
rect -6178 603178 -6006 603414
rect -6586 603094 -6006 603178
rect -6586 602858 -6414 603094
rect -6178 602858 -6006 603094
rect -6586 567414 -6006 602858
rect -6586 567178 -6414 567414
rect -6178 567178 -6006 567414
rect -6586 567094 -6006 567178
rect -6586 566858 -6414 567094
rect -6178 566858 -6006 567094
rect -6586 531414 -6006 566858
rect -6586 531178 -6414 531414
rect -6178 531178 -6006 531414
rect -6586 531094 -6006 531178
rect -6586 530858 -6414 531094
rect -6178 530858 -6006 531094
rect -6586 495414 -6006 530858
rect -6586 495178 -6414 495414
rect -6178 495178 -6006 495414
rect -6586 495094 -6006 495178
rect -6586 494858 -6414 495094
rect -6178 494858 -6006 495094
rect -6586 459414 -6006 494858
rect -6586 459178 -6414 459414
rect -6178 459178 -6006 459414
rect -6586 459094 -6006 459178
rect -6586 458858 -6414 459094
rect -6178 458858 -6006 459094
rect -6586 423414 -6006 458858
rect -6586 423178 -6414 423414
rect -6178 423178 -6006 423414
rect -6586 423094 -6006 423178
rect -6586 422858 -6414 423094
rect -6178 422858 -6006 423094
rect -6586 387414 -6006 422858
rect -6586 387178 -6414 387414
rect -6178 387178 -6006 387414
rect -6586 387094 -6006 387178
rect -6586 386858 -6414 387094
rect -6178 386858 -6006 387094
rect -6586 351414 -6006 386858
rect -6586 351178 -6414 351414
rect -6178 351178 -6006 351414
rect -6586 351094 -6006 351178
rect -6586 350858 -6414 351094
rect -6178 350858 -6006 351094
rect -6586 315414 -6006 350858
rect -6586 315178 -6414 315414
rect -6178 315178 -6006 315414
rect -6586 315094 -6006 315178
rect -6586 314858 -6414 315094
rect -6178 314858 -6006 315094
rect -6586 279414 -6006 314858
rect -6586 279178 -6414 279414
rect -6178 279178 -6006 279414
rect -6586 279094 -6006 279178
rect -6586 278858 -6414 279094
rect -6178 278858 -6006 279094
rect -6586 243414 -6006 278858
rect -6586 243178 -6414 243414
rect -6178 243178 -6006 243414
rect -6586 243094 -6006 243178
rect -6586 242858 -6414 243094
rect -6178 242858 -6006 243094
rect -6586 207414 -6006 242858
rect -6586 207178 -6414 207414
rect -6178 207178 -6006 207414
rect -6586 207094 -6006 207178
rect -6586 206858 -6414 207094
rect -6178 206858 -6006 207094
rect -6586 171414 -6006 206858
rect -6586 171178 -6414 171414
rect -6178 171178 -6006 171414
rect -6586 171094 -6006 171178
rect -6586 170858 -6414 171094
rect -6178 170858 -6006 171094
rect -6586 135414 -6006 170858
rect -6586 135178 -6414 135414
rect -6178 135178 -6006 135414
rect -6586 135094 -6006 135178
rect -6586 134858 -6414 135094
rect -6178 134858 -6006 135094
rect -6586 99414 -6006 134858
rect -6586 99178 -6414 99414
rect -6178 99178 -6006 99414
rect -6586 99094 -6006 99178
rect -6586 98858 -6414 99094
rect -6178 98858 -6006 99094
rect -6586 63414 -6006 98858
rect -6586 63178 -6414 63414
rect -6178 63178 -6006 63414
rect -6586 63094 -6006 63178
rect -6586 62858 -6414 63094
rect -6178 62858 -6006 63094
rect -6586 27414 -6006 62858
rect -6586 27178 -6414 27414
rect -6178 27178 -6006 27414
rect -6586 27094 -6006 27178
rect -6586 26858 -6414 27094
rect -6178 26858 -6006 27094
rect -6586 -4946 -6006 26858
rect -5666 708518 -5086 708530
rect -5666 708282 -5494 708518
rect -5258 708282 -5086 708518
rect -5666 708198 -5086 708282
rect -5666 707962 -5494 708198
rect -5258 707962 -5086 708198
rect -5666 693414 -5086 707962
rect 7774 708518 8354 709450
rect 7774 708282 7946 708518
rect 8182 708282 8354 708518
rect 7774 708198 8354 708282
rect 7774 707962 7946 708198
rect 8182 707962 8354 708198
rect -5666 693178 -5494 693414
rect -5258 693178 -5086 693414
rect -5666 693094 -5086 693178
rect -5666 692858 -5494 693094
rect -5258 692858 -5086 693094
rect -5666 657414 -5086 692858
rect -5666 657178 -5494 657414
rect -5258 657178 -5086 657414
rect -5666 657094 -5086 657178
rect -5666 656858 -5494 657094
rect -5258 656858 -5086 657094
rect -5666 621414 -5086 656858
rect -5666 621178 -5494 621414
rect -5258 621178 -5086 621414
rect -5666 621094 -5086 621178
rect -5666 620858 -5494 621094
rect -5258 620858 -5086 621094
rect -5666 585414 -5086 620858
rect -5666 585178 -5494 585414
rect -5258 585178 -5086 585414
rect -5666 585094 -5086 585178
rect -5666 584858 -5494 585094
rect -5258 584858 -5086 585094
rect -5666 549414 -5086 584858
rect -5666 549178 -5494 549414
rect -5258 549178 -5086 549414
rect -5666 549094 -5086 549178
rect -5666 548858 -5494 549094
rect -5258 548858 -5086 549094
rect -5666 513414 -5086 548858
rect -5666 513178 -5494 513414
rect -5258 513178 -5086 513414
rect -5666 513094 -5086 513178
rect -5666 512858 -5494 513094
rect -5258 512858 -5086 513094
rect -5666 477414 -5086 512858
rect -5666 477178 -5494 477414
rect -5258 477178 -5086 477414
rect -5666 477094 -5086 477178
rect -5666 476858 -5494 477094
rect -5258 476858 -5086 477094
rect -5666 441414 -5086 476858
rect -5666 441178 -5494 441414
rect -5258 441178 -5086 441414
rect -5666 441094 -5086 441178
rect -5666 440858 -5494 441094
rect -5258 440858 -5086 441094
rect -5666 405414 -5086 440858
rect -5666 405178 -5494 405414
rect -5258 405178 -5086 405414
rect -5666 405094 -5086 405178
rect -5666 404858 -5494 405094
rect -5258 404858 -5086 405094
rect -5666 369414 -5086 404858
rect -5666 369178 -5494 369414
rect -5258 369178 -5086 369414
rect -5666 369094 -5086 369178
rect -5666 368858 -5494 369094
rect -5258 368858 -5086 369094
rect -5666 333414 -5086 368858
rect -5666 333178 -5494 333414
rect -5258 333178 -5086 333414
rect -5666 333094 -5086 333178
rect -5666 332858 -5494 333094
rect -5258 332858 -5086 333094
rect -5666 297414 -5086 332858
rect -5666 297178 -5494 297414
rect -5258 297178 -5086 297414
rect -5666 297094 -5086 297178
rect -5666 296858 -5494 297094
rect -5258 296858 -5086 297094
rect -5666 261414 -5086 296858
rect -5666 261178 -5494 261414
rect -5258 261178 -5086 261414
rect -5666 261094 -5086 261178
rect -5666 260858 -5494 261094
rect -5258 260858 -5086 261094
rect -5666 225414 -5086 260858
rect -5666 225178 -5494 225414
rect -5258 225178 -5086 225414
rect -5666 225094 -5086 225178
rect -5666 224858 -5494 225094
rect -5258 224858 -5086 225094
rect -5666 189414 -5086 224858
rect -5666 189178 -5494 189414
rect -5258 189178 -5086 189414
rect -5666 189094 -5086 189178
rect -5666 188858 -5494 189094
rect -5258 188858 -5086 189094
rect -5666 153414 -5086 188858
rect -5666 153178 -5494 153414
rect -5258 153178 -5086 153414
rect -5666 153094 -5086 153178
rect -5666 152858 -5494 153094
rect -5258 152858 -5086 153094
rect -5666 117414 -5086 152858
rect -5666 117178 -5494 117414
rect -5258 117178 -5086 117414
rect -5666 117094 -5086 117178
rect -5666 116858 -5494 117094
rect -5258 116858 -5086 117094
rect -5666 81414 -5086 116858
rect -5666 81178 -5494 81414
rect -5258 81178 -5086 81414
rect -5666 81094 -5086 81178
rect -5666 80858 -5494 81094
rect -5258 80858 -5086 81094
rect -5666 45414 -5086 80858
rect -5666 45178 -5494 45414
rect -5258 45178 -5086 45414
rect -5666 45094 -5086 45178
rect -5666 44858 -5494 45094
rect -5258 44858 -5086 45094
rect -5666 9414 -5086 44858
rect -5666 9178 -5494 9414
rect -5258 9178 -5086 9414
rect -5666 9094 -5086 9178
rect -5666 8858 -5494 9094
rect -5258 8858 -5086 9094
rect -5666 -4026 -5086 8858
rect -4746 707598 -4166 707610
rect -4746 707362 -4574 707598
rect -4338 707362 -4166 707598
rect -4746 707278 -4166 707362
rect -4746 707042 -4574 707278
rect -4338 707042 -4166 707278
rect -4746 671934 -4166 707042
rect -4746 671698 -4574 671934
rect -4338 671698 -4166 671934
rect -4746 671614 -4166 671698
rect -4746 671378 -4574 671614
rect -4338 671378 -4166 671614
rect -4746 635934 -4166 671378
rect -4746 635698 -4574 635934
rect -4338 635698 -4166 635934
rect -4746 635614 -4166 635698
rect -4746 635378 -4574 635614
rect -4338 635378 -4166 635614
rect -4746 599934 -4166 635378
rect -4746 599698 -4574 599934
rect -4338 599698 -4166 599934
rect -4746 599614 -4166 599698
rect -4746 599378 -4574 599614
rect -4338 599378 -4166 599614
rect -4746 563934 -4166 599378
rect -4746 563698 -4574 563934
rect -4338 563698 -4166 563934
rect -4746 563614 -4166 563698
rect -4746 563378 -4574 563614
rect -4338 563378 -4166 563614
rect -4746 527934 -4166 563378
rect -4746 527698 -4574 527934
rect -4338 527698 -4166 527934
rect -4746 527614 -4166 527698
rect -4746 527378 -4574 527614
rect -4338 527378 -4166 527614
rect -4746 491934 -4166 527378
rect -4746 491698 -4574 491934
rect -4338 491698 -4166 491934
rect -4746 491614 -4166 491698
rect -4746 491378 -4574 491614
rect -4338 491378 -4166 491614
rect -4746 455934 -4166 491378
rect -4746 455698 -4574 455934
rect -4338 455698 -4166 455934
rect -4746 455614 -4166 455698
rect -4746 455378 -4574 455614
rect -4338 455378 -4166 455614
rect -4746 419934 -4166 455378
rect -4746 419698 -4574 419934
rect -4338 419698 -4166 419934
rect -4746 419614 -4166 419698
rect -4746 419378 -4574 419614
rect -4338 419378 -4166 419614
rect -4746 383934 -4166 419378
rect -4746 383698 -4574 383934
rect -4338 383698 -4166 383934
rect -4746 383614 -4166 383698
rect -4746 383378 -4574 383614
rect -4338 383378 -4166 383614
rect -4746 347934 -4166 383378
rect -4746 347698 -4574 347934
rect -4338 347698 -4166 347934
rect -4746 347614 -4166 347698
rect -4746 347378 -4574 347614
rect -4338 347378 -4166 347614
rect -4746 311934 -4166 347378
rect -4746 311698 -4574 311934
rect -4338 311698 -4166 311934
rect -4746 311614 -4166 311698
rect -4746 311378 -4574 311614
rect -4338 311378 -4166 311614
rect -4746 275934 -4166 311378
rect -4746 275698 -4574 275934
rect -4338 275698 -4166 275934
rect -4746 275614 -4166 275698
rect -4746 275378 -4574 275614
rect -4338 275378 -4166 275614
rect -4746 239934 -4166 275378
rect -4746 239698 -4574 239934
rect -4338 239698 -4166 239934
rect -4746 239614 -4166 239698
rect -4746 239378 -4574 239614
rect -4338 239378 -4166 239614
rect -4746 203934 -4166 239378
rect -4746 203698 -4574 203934
rect -4338 203698 -4166 203934
rect -4746 203614 -4166 203698
rect -4746 203378 -4574 203614
rect -4338 203378 -4166 203614
rect -4746 167934 -4166 203378
rect -4746 167698 -4574 167934
rect -4338 167698 -4166 167934
rect -4746 167614 -4166 167698
rect -4746 167378 -4574 167614
rect -4338 167378 -4166 167614
rect -4746 131934 -4166 167378
rect -4746 131698 -4574 131934
rect -4338 131698 -4166 131934
rect -4746 131614 -4166 131698
rect -4746 131378 -4574 131614
rect -4338 131378 -4166 131614
rect -4746 95934 -4166 131378
rect -4746 95698 -4574 95934
rect -4338 95698 -4166 95934
rect -4746 95614 -4166 95698
rect -4746 95378 -4574 95614
rect -4338 95378 -4166 95614
rect -4746 59934 -4166 95378
rect -4746 59698 -4574 59934
rect -4338 59698 -4166 59934
rect -4746 59614 -4166 59698
rect -4746 59378 -4574 59614
rect -4338 59378 -4166 59614
rect -4746 23934 -4166 59378
rect -4746 23698 -4574 23934
rect -4338 23698 -4166 23934
rect -4746 23614 -4166 23698
rect -4746 23378 -4574 23614
rect -4338 23378 -4166 23614
rect -4746 -3106 -4166 23378
rect -3826 706678 -3246 706690
rect -3826 706442 -3654 706678
rect -3418 706442 -3246 706678
rect -3826 706358 -3246 706442
rect -3826 706122 -3654 706358
rect -3418 706122 -3246 706358
rect -3826 689934 -3246 706122
rect 4294 706678 4874 707610
rect 4294 706442 4466 706678
rect 4702 706442 4874 706678
rect 4294 706358 4874 706442
rect 4294 706122 4466 706358
rect 4702 706122 4874 706358
rect -3826 689698 -3654 689934
rect -3418 689698 -3246 689934
rect -3826 689614 -3246 689698
rect -3826 689378 -3654 689614
rect -3418 689378 -3246 689614
rect -3826 653934 -3246 689378
rect -3826 653698 -3654 653934
rect -3418 653698 -3246 653934
rect -3826 653614 -3246 653698
rect -3826 653378 -3654 653614
rect -3418 653378 -3246 653614
rect -3826 617934 -3246 653378
rect -3826 617698 -3654 617934
rect -3418 617698 -3246 617934
rect -3826 617614 -3246 617698
rect -3826 617378 -3654 617614
rect -3418 617378 -3246 617614
rect -3826 581934 -3246 617378
rect -3826 581698 -3654 581934
rect -3418 581698 -3246 581934
rect -3826 581614 -3246 581698
rect -3826 581378 -3654 581614
rect -3418 581378 -3246 581614
rect -3826 545934 -3246 581378
rect -3826 545698 -3654 545934
rect -3418 545698 -3246 545934
rect -3826 545614 -3246 545698
rect -3826 545378 -3654 545614
rect -3418 545378 -3246 545614
rect -3826 509934 -3246 545378
rect -3826 509698 -3654 509934
rect -3418 509698 -3246 509934
rect -3826 509614 -3246 509698
rect -3826 509378 -3654 509614
rect -3418 509378 -3246 509614
rect -3826 473934 -3246 509378
rect -3826 473698 -3654 473934
rect -3418 473698 -3246 473934
rect -3826 473614 -3246 473698
rect -3826 473378 -3654 473614
rect -3418 473378 -3246 473614
rect -3826 437934 -3246 473378
rect -3826 437698 -3654 437934
rect -3418 437698 -3246 437934
rect -3826 437614 -3246 437698
rect -3826 437378 -3654 437614
rect -3418 437378 -3246 437614
rect -3826 401934 -3246 437378
rect -3826 401698 -3654 401934
rect -3418 401698 -3246 401934
rect -3826 401614 -3246 401698
rect -3826 401378 -3654 401614
rect -3418 401378 -3246 401614
rect -3826 365934 -3246 401378
rect -3826 365698 -3654 365934
rect -3418 365698 -3246 365934
rect -3826 365614 -3246 365698
rect -3826 365378 -3654 365614
rect -3418 365378 -3246 365614
rect -3826 329934 -3246 365378
rect -3826 329698 -3654 329934
rect -3418 329698 -3246 329934
rect -3826 329614 -3246 329698
rect -3826 329378 -3654 329614
rect -3418 329378 -3246 329614
rect -3826 293934 -3246 329378
rect -3826 293698 -3654 293934
rect -3418 293698 -3246 293934
rect -3826 293614 -3246 293698
rect -3826 293378 -3654 293614
rect -3418 293378 -3246 293614
rect -3826 257934 -3246 293378
rect -3826 257698 -3654 257934
rect -3418 257698 -3246 257934
rect -3826 257614 -3246 257698
rect -3826 257378 -3654 257614
rect -3418 257378 -3246 257614
rect -3826 221934 -3246 257378
rect -3826 221698 -3654 221934
rect -3418 221698 -3246 221934
rect -3826 221614 -3246 221698
rect -3826 221378 -3654 221614
rect -3418 221378 -3246 221614
rect -3826 185934 -3246 221378
rect -3826 185698 -3654 185934
rect -3418 185698 -3246 185934
rect -3826 185614 -3246 185698
rect -3826 185378 -3654 185614
rect -3418 185378 -3246 185614
rect -3826 149934 -3246 185378
rect -3826 149698 -3654 149934
rect -3418 149698 -3246 149934
rect -3826 149614 -3246 149698
rect -3826 149378 -3654 149614
rect -3418 149378 -3246 149614
rect -3826 113934 -3246 149378
rect -3826 113698 -3654 113934
rect -3418 113698 -3246 113934
rect -3826 113614 -3246 113698
rect -3826 113378 -3654 113614
rect -3418 113378 -3246 113614
rect -3826 77934 -3246 113378
rect -3826 77698 -3654 77934
rect -3418 77698 -3246 77934
rect -3826 77614 -3246 77698
rect -3826 77378 -3654 77614
rect -3418 77378 -3246 77614
rect -3826 41934 -3246 77378
rect -3826 41698 -3654 41934
rect -3418 41698 -3246 41934
rect -3826 41614 -3246 41698
rect -3826 41378 -3654 41614
rect -3418 41378 -3246 41614
rect -3826 5934 -3246 41378
rect -3826 5698 -3654 5934
rect -3418 5698 -3246 5934
rect -3826 5614 -3246 5698
rect -3826 5378 -3654 5614
rect -3418 5378 -3246 5614
rect -3826 -2186 -3246 5378
rect -2906 705758 -2326 705770
rect -2906 705522 -2734 705758
rect -2498 705522 -2326 705758
rect -2906 705438 -2326 705522
rect -2906 705202 -2734 705438
rect -2498 705202 -2326 705438
rect -2906 668454 -2326 705202
rect -2906 668218 -2734 668454
rect -2498 668218 -2326 668454
rect -2906 668134 -2326 668218
rect -2906 667898 -2734 668134
rect -2498 667898 -2326 668134
rect -2906 632454 -2326 667898
rect -2906 632218 -2734 632454
rect -2498 632218 -2326 632454
rect -2906 632134 -2326 632218
rect -2906 631898 -2734 632134
rect -2498 631898 -2326 632134
rect -2906 596454 -2326 631898
rect -2906 596218 -2734 596454
rect -2498 596218 -2326 596454
rect -2906 596134 -2326 596218
rect -2906 595898 -2734 596134
rect -2498 595898 -2326 596134
rect -2906 560454 -2326 595898
rect -2906 560218 -2734 560454
rect -2498 560218 -2326 560454
rect -2906 560134 -2326 560218
rect -2906 559898 -2734 560134
rect -2498 559898 -2326 560134
rect -2906 524454 -2326 559898
rect -2906 524218 -2734 524454
rect -2498 524218 -2326 524454
rect -2906 524134 -2326 524218
rect -2906 523898 -2734 524134
rect -2498 523898 -2326 524134
rect -2906 488454 -2326 523898
rect -2906 488218 -2734 488454
rect -2498 488218 -2326 488454
rect -2906 488134 -2326 488218
rect -2906 487898 -2734 488134
rect -2498 487898 -2326 488134
rect -2906 452454 -2326 487898
rect -2906 452218 -2734 452454
rect -2498 452218 -2326 452454
rect -2906 452134 -2326 452218
rect -2906 451898 -2734 452134
rect -2498 451898 -2326 452134
rect -2906 416454 -2326 451898
rect -2906 416218 -2734 416454
rect -2498 416218 -2326 416454
rect -2906 416134 -2326 416218
rect -2906 415898 -2734 416134
rect -2498 415898 -2326 416134
rect -2906 380454 -2326 415898
rect -2906 380218 -2734 380454
rect -2498 380218 -2326 380454
rect -2906 380134 -2326 380218
rect -2906 379898 -2734 380134
rect -2498 379898 -2326 380134
rect -2906 344454 -2326 379898
rect -2906 344218 -2734 344454
rect -2498 344218 -2326 344454
rect -2906 344134 -2326 344218
rect -2906 343898 -2734 344134
rect -2498 343898 -2326 344134
rect -2906 308454 -2326 343898
rect -2906 308218 -2734 308454
rect -2498 308218 -2326 308454
rect -2906 308134 -2326 308218
rect -2906 307898 -2734 308134
rect -2498 307898 -2326 308134
rect -2906 272454 -2326 307898
rect -2906 272218 -2734 272454
rect -2498 272218 -2326 272454
rect -2906 272134 -2326 272218
rect -2906 271898 -2734 272134
rect -2498 271898 -2326 272134
rect -2906 236454 -2326 271898
rect -2906 236218 -2734 236454
rect -2498 236218 -2326 236454
rect -2906 236134 -2326 236218
rect -2906 235898 -2734 236134
rect -2498 235898 -2326 236134
rect -2906 200454 -2326 235898
rect -2906 200218 -2734 200454
rect -2498 200218 -2326 200454
rect -2906 200134 -2326 200218
rect -2906 199898 -2734 200134
rect -2498 199898 -2326 200134
rect -2906 164454 -2326 199898
rect -2906 164218 -2734 164454
rect -2498 164218 -2326 164454
rect -2906 164134 -2326 164218
rect -2906 163898 -2734 164134
rect -2498 163898 -2326 164134
rect -2906 128454 -2326 163898
rect -2906 128218 -2734 128454
rect -2498 128218 -2326 128454
rect -2906 128134 -2326 128218
rect -2906 127898 -2734 128134
rect -2498 127898 -2326 128134
rect -2906 92454 -2326 127898
rect -2906 92218 -2734 92454
rect -2498 92218 -2326 92454
rect -2906 92134 -2326 92218
rect -2906 91898 -2734 92134
rect -2498 91898 -2326 92134
rect -2906 56454 -2326 91898
rect -2906 56218 -2734 56454
rect -2498 56218 -2326 56454
rect -2906 56134 -2326 56218
rect -2906 55898 -2734 56134
rect -2498 55898 -2326 56134
rect -2906 20454 -2326 55898
rect -2906 20218 -2734 20454
rect -2498 20218 -2326 20454
rect -2906 20134 -2326 20218
rect -2906 19898 -2734 20134
rect -2498 19898 -2326 20134
rect -2906 -1266 -2326 19898
rect -1986 704838 -1406 704850
rect -1986 704602 -1814 704838
rect -1578 704602 -1406 704838
rect -1986 704518 -1406 704602
rect -1986 704282 -1814 704518
rect -1578 704282 -1406 704518
rect -1986 686454 -1406 704282
rect -1986 686218 -1814 686454
rect -1578 686218 -1406 686454
rect -1986 686134 -1406 686218
rect -1986 685898 -1814 686134
rect -1578 685898 -1406 686134
rect -1986 650454 -1406 685898
rect -1986 650218 -1814 650454
rect -1578 650218 -1406 650454
rect -1986 650134 -1406 650218
rect -1986 649898 -1814 650134
rect -1578 649898 -1406 650134
rect -1986 614454 -1406 649898
rect -1986 614218 -1814 614454
rect -1578 614218 -1406 614454
rect -1986 614134 -1406 614218
rect -1986 613898 -1814 614134
rect -1578 613898 -1406 614134
rect -1986 578454 -1406 613898
rect -1986 578218 -1814 578454
rect -1578 578218 -1406 578454
rect -1986 578134 -1406 578218
rect -1986 577898 -1814 578134
rect -1578 577898 -1406 578134
rect -1986 542454 -1406 577898
rect -1986 542218 -1814 542454
rect -1578 542218 -1406 542454
rect -1986 542134 -1406 542218
rect -1986 541898 -1814 542134
rect -1578 541898 -1406 542134
rect -1986 506454 -1406 541898
rect -1986 506218 -1814 506454
rect -1578 506218 -1406 506454
rect -1986 506134 -1406 506218
rect -1986 505898 -1814 506134
rect -1578 505898 -1406 506134
rect -1986 470454 -1406 505898
rect -1986 470218 -1814 470454
rect -1578 470218 -1406 470454
rect -1986 470134 -1406 470218
rect -1986 469898 -1814 470134
rect -1578 469898 -1406 470134
rect -1986 434454 -1406 469898
rect -1986 434218 -1814 434454
rect -1578 434218 -1406 434454
rect -1986 434134 -1406 434218
rect -1986 433898 -1814 434134
rect -1578 433898 -1406 434134
rect -1986 398454 -1406 433898
rect -1986 398218 -1814 398454
rect -1578 398218 -1406 398454
rect -1986 398134 -1406 398218
rect -1986 397898 -1814 398134
rect -1578 397898 -1406 398134
rect -1986 362454 -1406 397898
rect -1986 362218 -1814 362454
rect -1578 362218 -1406 362454
rect -1986 362134 -1406 362218
rect -1986 361898 -1814 362134
rect -1578 361898 -1406 362134
rect -1986 326454 -1406 361898
rect -1986 326218 -1814 326454
rect -1578 326218 -1406 326454
rect -1986 326134 -1406 326218
rect -1986 325898 -1814 326134
rect -1578 325898 -1406 326134
rect -1986 290454 -1406 325898
rect -1986 290218 -1814 290454
rect -1578 290218 -1406 290454
rect -1986 290134 -1406 290218
rect -1986 289898 -1814 290134
rect -1578 289898 -1406 290134
rect -1986 254454 -1406 289898
rect -1986 254218 -1814 254454
rect -1578 254218 -1406 254454
rect -1986 254134 -1406 254218
rect -1986 253898 -1814 254134
rect -1578 253898 -1406 254134
rect -1986 218454 -1406 253898
rect -1986 218218 -1814 218454
rect -1578 218218 -1406 218454
rect -1986 218134 -1406 218218
rect -1986 217898 -1814 218134
rect -1578 217898 -1406 218134
rect -1986 182454 -1406 217898
rect -1986 182218 -1814 182454
rect -1578 182218 -1406 182454
rect -1986 182134 -1406 182218
rect -1986 181898 -1814 182134
rect -1578 181898 -1406 182134
rect -1986 146454 -1406 181898
rect -1986 146218 -1814 146454
rect -1578 146218 -1406 146454
rect -1986 146134 -1406 146218
rect -1986 145898 -1814 146134
rect -1578 145898 -1406 146134
rect -1986 110454 -1406 145898
rect -1986 110218 -1814 110454
rect -1578 110218 -1406 110454
rect -1986 110134 -1406 110218
rect -1986 109898 -1814 110134
rect -1578 109898 -1406 110134
rect -1986 74454 -1406 109898
rect -1986 74218 -1814 74454
rect -1578 74218 -1406 74454
rect -1986 74134 -1406 74218
rect -1986 73898 -1814 74134
rect -1578 73898 -1406 74134
rect -1986 38454 -1406 73898
rect -1986 38218 -1814 38454
rect -1578 38218 -1406 38454
rect -1986 38134 -1406 38218
rect -1986 37898 -1814 38134
rect -1578 37898 -1406 38134
rect -1986 2454 -1406 37898
rect -1986 2218 -1814 2454
rect -1578 2218 -1406 2454
rect -1986 2134 -1406 2218
rect -1986 1898 -1814 2134
rect -1578 1898 -1406 2134
rect -1986 -346 -1406 1898
rect -1986 -582 -1814 -346
rect -1578 -582 -1406 -346
rect -1986 -666 -1406 -582
rect -1986 -902 -1814 -666
rect -1578 -902 -1406 -666
rect -1986 -914 -1406 -902
rect 814 704838 1394 705770
rect 814 704602 986 704838
rect 1222 704602 1394 704838
rect 814 704518 1394 704602
rect 814 704282 986 704518
rect 1222 704282 1394 704518
rect 814 686454 1394 704282
rect 814 686218 986 686454
rect 1222 686218 1394 686454
rect 814 686134 1394 686218
rect 814 685898 986 686134
rect 1222 685898 1394 686134
rect 814 650454 1394 685898
rect 814 650218 986 650454
rect 1222 650218 1394 650454
rect 814 650134 1394 650218
rect 814 649898 986 650134
rect 1222 649898 1394 650134
rect 814 614454 1394 649898
rect 814 614218 986 614454
rect 1222 614218 1394 614454
rect 814 614134 1394 614218
rect 814 613898 986 614134
rect 1222 613898 1394 614134
rect 814 578454 1394 613898
rect 814 578218 986 578454
rect 1222 578218 1394 578454
rect 814 578134 1394 578218
rect 814 577898 986 578134
rect 1222 577898 1394 578134
rect 814 542454 1394 577898
rect 814 542218 986 542454
rect 1222 542218 1394 542454
rect 814 542134 1394 542218
rect 814 541898 986 542134
rect 1222 541898 1394 542134
rect 814 506454 1394 541898
rect 814 506218 986 506454
rect 1222 506218 1394 506454
rect 814 506134 1394 506218
rect 814 505898 986 506134
rect 1222 505898 1394 506134
rect 814 470454 1394 505898
rect 814 470218 986 470454
rect 1222 470218 1394 470454
rect 814 470134 1394 470218
rect 814 469898 986 470134
rect 1222 469898 1394 470134
rect 814 434454 1394 469898
rect 814 434218 986 434454
rect 1222 434218 1394 434454
rect 814 434134 1394 434218
rect 814 433898 986 434134
rect 1222 433898 1394 434134
rect 814 398454 1394 433898
rect 814 398218 986 398454
rect 1222 398218 1394 398454
rect 814 398134 1394 398218
rect 814 397898 986 398134
rect 1222 397898 1394 398134
rect 814 362454 1394 397898
rect 814 362218 986 362454
rect 1222 362218 1394 362454
rect 814 362134 1394 362218
rect 814 361898 986 362134
rect 1222 361898 1394 362134
rect 814 326454 1394 361898
rect 814 326218 986 326454
rect 1222 326218 1394 326454
rect 814 326134 1394 326218
rect 814 325898 986 326134
rect 1222 325898 1394 326134
rect 814 290454 1394 325898
rect 814 290218 986 290454
rect 1222 290218 1394 290454
rect 814 290134 1394 290218
rect 814 289898 986 290134
rect 1222 289898 1394 290134
rect 814 254454 1394 289898
rect 814 254218 986 254454
rect 1222 254218 1394 254454
rect 814 254134 1394 254218
rect 814 253898 986 254134
rect 1222 253898 1394 254134
rect 814 218454 1394 253898
rect 814 218218 986 218454
rect 1222 218218 1394 218454
rect 814 218134 1394 218218
rect 814 217898 986 218134
rect 1222 217898 1394 218134
rect 814 182454 1394 217898
rect 814 182218 986 182454
rect 1222 182218 1394 182454
rect 814 182134 1394 182218
rect 814 181898 986 182134
rect 1222 181898 1394 182134
rect 814 146454 1394 181898
rect 814 146218 986 146454
rect 1222 146218 1394 146454
rect 814 146134 1394 146218
rect 814 145898 986 146134
rect 1222 145898 1394 146134
rect 814 110454 1394 145898
rect 814 110218 986 110454
rect 1222 110218 1394 110454
rect 814 110134 1394 110218
rect 814 109898 986 110134
rect 1222 109898 1394 110134
rect 814 74454 1394 109898
rect 814 74218 986 74454
rect 1222 74218 1394 74454
rect 814 74134 1394 74218
rect 814 73898 986 74134
rect 1222 73898 1394 74134
rect 814 38454 1394 73898
rect 814 38218 986 38454
rect 1222 38218 1394 38454
rect 814 38134 1394 38218
rect 814 37898 986 38134
rect 1222 37898 1394 38134
rect 814 2454 1394 37898
rect 814 2218 986 2454
rect 1222 2218 1394 2454
rect 814 2134 1394 2218
rect 814 1898 986 2134
rect 1222 1898 1394 2134
rect 814 -346 1394 1898
rect 814 -582 986 -346
rect 1222 -582 1394 -346
rect 814 -666 1394 -582
rect 814 -902 986 -666
rect 1222 -902 1394 -666
rect -2906 -1502 -2734 -1266
rect -2498 -1502 -2326 -1266
rect -2906 -1586 -2326 -1502
rect -2906 -1822 -2734 -1586
rect -2498 -1822 -2326 -1586
rect -2906 -1834 -2326 -1822
rect 814 -1834 1394 -902
rect 4294 689934 4874 706122
rect 4294 689698 4466 689934
rect 4702 689698 4874 689934
rect 4294 689614 4874 689698
rect 4294 689378 4466 689614
rect 4702 689378 4874 689614
rect 4294 653934 4874 689378
rect 4294 653698 4466 653934
rect 4702 653698 4874 653934
rect 4294 653614 4874 653698
rect 4294 653378 4466 653614
rect 4702 653378 4874 653614
rect 4294 617934 4874 653378
rect 4294 617698 4466 617934
rect 4702 617698 4874 617934
rect 4294 617614 4874 617698
rect 4294 617378 4466 617614
rect 4702 617378 4874 617614
rect 4294 581934 4874 617378
rect 4294 581698 4466 581934
rect 4702 581698 4874 581934
rect 4294 581614 4874 581698
rect 4294 581378 4466 581614
rect 4702 581378 4874 581614
rect 4294 545934 4874 581378
rect 4294 545698 4466 545934
rect 4702 545698 4874 545934
rect 4294 545614 4874 545698
rect 4294 545378 4466 545614
rect 4702 545378 4874 545614
rect 4294 509934 4874 545378
rect 4294 509698 4466 509934
rect 4702 509698 4874 509934
rect 4294 509614 4874 509698
rect 4294 509378 4466 509614
rect 4702 509378 4874 509614
rect 4294 473934 4874 509378
rect 4294 473698 4466 473934
rect 4702 473698 4874 473934
rect 4294 473614 4874 473698
rect 4294 473378 4466 473614
rect 4702 473378 4874 473614
rect 4294 437934 4874 473378
rect 4294 437698 4466 437934
rect 4702 437698 4874 437934
rect 4294 437614 4874 437698
rect 4294 437378 4466 437614
rect 4702 437378 4874 437614
rect 4294 401934 4874 437378
rect 4294 401698 4466 401934
rect 4702 401698 4874 401934
rect 4294 401614 4874 401698
rect 4294 401378 4466 401614
rect 4702 401378 4874 401614
rect 4294 365934 4874 401378
rect 4294 365698 4466 365934
rect 4702 365698 4874 365934
rect 4294 365614 4874 365698
rect 4294 365378 4466 365614
rect 4702 365378 4874 365614
rect 4294 329934 4874 365378
rect 4294 329698 4466 329934
rect 4702 329698 4874 329934
rect 4294 329614 4874 329698
rect 4294 329378 4466 329614
rect 4702 329378 4874 329614
rect 4294 293934 4874 329378
rect 4294 293698 4466 293934
rect 4702 293698 4874 293934
rect 4294 293614 4874 293698
rect 4294 293378 4466 293614
rect 4702 293378 4874 293614
rect 4294 257934 4874 293378
rect 4294 257698 4466 257934
rect 4702 257698 4874 257934
rect 4294 257614 4874 257698
rect 4294 257378 4466 257614
rect 4702 257378 4874 257614
rect 4294 221934 4874 257378
rect 4294 221698 4466 221934
rect 4702 221698 4874 221934
rect 4294 221614 4874 221698
rect 4294 221378 4466 221614
rect 4702 221378 4874 221614
rect 4294 185934 4874 221378
rect 4294 185698 4466 185934
rect 4702 185698 4874 185934
rect 4294 185614 4874 185698
rect 4294 185378 4466 185614
rect 4702 185378 4874 185614
rect 4294 149934 4874 185378
rect 4294 149698 4466 149934
rect 4702 149698 4874 149934
rect 4294 149614 4874 149698
rect 4294 149378 4466 149614
rect 4702 149378 4874 149614
rect 4294 113934 4874 149378
rect 4294 113698 4466 113934
rect 4702 113698 4874 113934
rect 4294 113614 4874 113698
rect 4294 113378 4466 113614
rect 4702 113378 4874 113614
rect 4294 77934 4874 113378
rect 4294 77698 4466 77934
rect 4702 77698 4874 77934
rect 4294 77614 4874 77698
rect 4294 77378 4466 77614
rect 4702 77378 4874 77614
rect 4294 41934 4874 77378
rect 4294 41698 4466 41934
rect 4702 41698 4874 41934
rect 4294 41614 4874 41698
rect 4294 41378 4466 41614
rect 4702 41378 4874 41614
rect 4294 5934 4874 41378
rect 4294 5698 4466 5934
rect 4702 5698 4874 5934
rect 4294 5614 4874 5698
rect 4294 5378 4466 5614
rect 4702 5378 4874 5614
rect -3826 -2422 -3654 -2186
rect -3418 -2422 -3246 -2186
rect -3826 -2506 -3246 -2422
rect -3826 -2742 -3654 -2506
rect -3418 -2742 -3246 -2506
rect -3826 -2754 -3246 -2742
rect 4294 -2186 4874 5378
rect 4294 -2422 4466 -2186
rect 4702 -2422 4874 -2186
rect 4294 -2506 4874 -2422
rect 4294 -2742 4466 -2506
rect 4702 -2742 4874 -2506
rect -4746 -3342 -4574 -3106
rect -4338 -3342 -4166 -3106
rect -4746 -3426 -4166 -3342
rect -4746 -3662 -4574 -3426
rect -4338 -3662 -4166 -3426
rect -4746 -3674 -4166 -3662
rect 4294 -3674 4874 -2742
rect 7774 693414 8354 707962
rect 7774 693178 7946 693414
rect 8182 693178 8354 693414
rect 7774 693094 8354 693178
rect 7774 692858 7946 693094
rect 8182 692858 8354 693094
rect 7774 657414 8354 692858
rect 7774 657178 7946 657414
rect 8182 657178 8354 657414
rect 7774 657094 8354 657178
rect 7774 656858 7946 657094
rect 8182 656858 8354 657094
rect 7774 621414 8354 656858
rect 7774 621178 7946 621414
rect 8182 621178 8354 621414
rect 7774 621094 8354 621178
rect 7774 620858 7946 621094
rect 8182 620858 8354 621094
rect 7774 585414 8354 620858
rect 7774 585178 7946 585414
rect 8182 585178 8354 585414
rect 7774 585094 8354 585178
rect 7774 584858 7946 585094
rect 8182 584858 8354 585094
rect 7774 549414 8354 584858
rect 7774 549178 7946 549414
rect 8182 549178 8354 549414
rect 7774 549094 8354 549178
rect 7774 548858 7946 549094
rect 8182 548858 8354 549094
rect 7774 513414 8354 548858
rect 7774 513178 7946 513414
rect 8182 513178 8354 513414
rect 7774 513094 8354 513178
rect 7774 512858 7946 513094
rect 8182 512858 8354 513094
rect 7774 477414 8354 512858
rect 7774 477178 7946 477414
rect 8182 477178 8354 477414
rect 7774 477094 8354 477178
rect 7774 476858 7946 477094
rect 8182 476858 8354 477094
rect 7774 441414 8354 476858
rect 7774 441178 7946 441414
rect 8182 441178 8354 441414
rect 7774 441094 8354 441178
rect 7774 440858 7946 441094
rect 8182 440858 8354 441094
rect 7774 405414 8354 440858
rect 7774 405178 7946 405414
rect 8182 405178 8354 405414
rect 7774 405094 8354 405178
rect 7774 404858 7946 405094
rect 8182 404858 8354 405094
rect 7774 369414 8354 404858
rect 7774 369178 7946 369414
rect 8182 369178 8354 369414
rect 7774 369094 8354 369178
rect 7774 368858 7946 369094
rect 8182 368858 8354 369094
rect 7774 333414 8354 368858
rect 7774 333178 7946 333414
rect 8182 333178 8354 333414
rect 7774 333094 8354 333178
rect 7774 332858 7946 333094
rect 8182 332858 8354 333094
rect 7774 297414 8354 332858
rect 7774 297178 7946 297414
rect 8182 297178 8354 297414
rect 7774 297094 8354 297178
rect 7774 296858 7946 297094
rect 8182 296858 8354 297094
rect 7774 261414 8354 296858
rect 7774 261178 7946 261414
rect 8182 261178 8354 261414
rect 7774 261094 8354 261178
rect 7774 260858 7946 261094
rect 8182 260858 8354 261094
rect 7774 225414 8354 260858
rect 7774 225178 7946 225414
rect 8182 225178 8354 225414
rect 7774 225094 8354 225178
rect 7774 224858 7946 225094
rect 8182 224858 8354 225094
rect 7774 189414 8354 224858
rect 7774 189178 7946 189414
rect 8182 189178 8354 189414
rect 7774 189094 8354 189178
rect 7774 188858 7946 189094
rect 8182 188858 8354 189094
rect 7774 153414 8354 188858
rect 7774 153178 7946 153414
rect 8182 153178 8354 153414
rect 7774 153094 8354 153178
rect 7774 152858 7946 153094
rect 8182 152858 8354 153094
rect 7774 117414 8354 152858
rect 7774 117178 7946 117414
rect 8182 117178 8354 117414
rect 7774 117094 8354 117178
rect 7774 116858 7946 117094
rect 8182 116858 8354 117094
rect 7774 81414 8354 116858
rect 7774 81178 7946 81414
rect 8182 81178 8354 81414
rect 7774 81094 8354 81178
rect 7774 80858 7946 81094
rect 8182 80858 8354 81094
rect 7774 45414 8354 80858
rect 7774 45178 7946 45414
rect 8182 45178 8354 45414
rect 7774 45094 8354 45178
rect 7774 44858 7946 45094
rect 8182 44858 8354 45094
rect 7774 9414 8354 44858
rect 7774 9178 7946 9414
rect 8182 9178 8354 9414
rect 7774 9094 8354 9178
rect 7774 8858 7946 9094
rect 8182 8858 8354 9094
rect -5666 -4262 -5494 -4026
rect -5258 -4262 -5086 -4026
rect -5666 -4346 -5086 -4262
rect -5666 -4582 -5494 -4346
rect -5258 -4582 -5086 -4346
rect -5666 -4594 -5086 -4582
rect 7774 -4026 8354 8858
rect 7774 -4262 7946 -4026
rect 8182 -4262 8354 -4026
rect 7774 -4346 8354 -4262
rect 7774 -4582 7946 -4346
rect 8182 -4582 8354 -4346
rect -6586 -5182 -6414 -4946
rect -6178 -5182 -6006 -4946
rect -6586 -5266 -6006 -5182
rect -6586 -5502 -6414 -5266
rect -6178 -5502 -6006 -5266
rect -6586 -5514 -6006 -5502
rect 7774 -5514 8354 -4582
rect 11254 696894 11834 709802
rect 29254 711278 29834 711290
rect 29254 711042 29426 711278
rect 29662 711042 29834 711278
rect 29254 710958 29834 711042
rect 29254 710722 29426 710958
rect 29662 710722 29834 710958
rect 25774 709438 26354 709450
rect 25774 709202 25946 709438
rect 26182 709202 26354 709438
rect 25774 709118 26354 709202
rect 25774 708882 25946 709118
rect 26182 708882 26354 709118
rect 22294 707598 22874 707610
rect 22294 707362 22466 707598
rect 22702 707362 22874 707598
rect 22294 707278 22874 707362
rect 22294 707042 22466 707278
rect 22702 707042 22874 707278
rect 11254 696658 11426 696894
rect 11662 696658 11834 696894
rect 11254 696574 11834 696658
rect 11254 696338 11426 696574
rect 11662 696338 11834 696574
rect 11254 660894 11834 696338
rect 11254 660658 11426 660894
rect 11662 660658 11834 660894
rect 11254 660574 11834 660658
rect 11254 660338 11426 660574
rect 11662 660338 11834 660574
rect 11254 624894 11834 660338
rect 11254 624658 11426 624894
rect 11662 624658 11834 624894
rect 11254 624574 11834 624658
rect 11254 624338 11426 624574
rect 11662 624338 11834 624574
rect 11254 588894 11834 624338
rect 11254 588658 11426 588894
rect 11662 588658 11834 588894
rect 11254 588574 11834 588658
rect 11254 588338 11426 588574
rect 11662 588338 11834 588574
rect 11254 552894 11834 588338
rect 11254 552658 11426 552894
rect 11662 552658 11834 552894
rect 11254 552574 11834 552658
rect 11254 552338 11426 552574
rect 11662 552338 11834 552574
rect 11254 516894 11834 552338
rect 11254 516658 11426 516894
rect 11662 516658 11834 516894
rect 11254 516574 11834 516658
rect 11254 516338 11426 516574
rect 11662 516338 11834 516574
rect 11254 480894 11834 516338
rect 11254 480658 11426 480894
rect 11662 480658 11834 480894
rect 11254 480574 11834 480658
rect 11254 480338 11426 480574
rect 11662 480338 11834 480574
rect 11254 444894 11834 480338
rect 11254 444658 11426 444894
rect 11662 444658 11834 444894
rect 11254 444574 11834 444658
rect 11254 444338 11426 444574
rect 11662 444338 11834 444574
rect 11254 408894 11834 444338
rect 11254 408658 11426 408894
rect 11662 408658 11834 408894
rect 11254 408574 11834 408658
rect 11254 408338 11426 408574
rect 11662 408338 11834 408574
rect 11254 372894 11834 408338
rect 11254 372658 11426 372894
rect 11662 372658 11834 372894
rect 11254 372574 11834 372658
rect 11254 372338 11426 372574
rect 11662 372338 11834 372574
rect 11254 336894 11834 372338
rect 11254 336658 11426 336894
rect 11662 336658 11834 336894
rect 11254 336574 11834 336658
rect 11254 336338 11426 336574
rect 11662 336338 11834 336574
rect 11254 300894 11834 336338
rect 11254 300658 11426 300894
rect 11662 300658 11834 300894
rect 11254 300574 11834 300658
rect 11254 300338 11426 300574
rect 11662 300338 11834 300574
rect 11254 264894 11834 300338
rect 11254 264658 11426 264894
rect 11662 264658 11834 264894
rect 11254 264574 11834 264658
rect 11254 264338 11426 264574
rect 11662 264338 11834 264574
rect 11254 228894 11834 264338
rect 11254 228658 11426 228894
rect 11662 228658 11834 228894
rect 11254 228574 11834 228658
rect 11254 228338 11426 228574
rect 11662 228338 11834 228574
rect 11254 192894 11834 228338
rect 11254 192658 11426 192894
rect 11662 192658 11834 192894
rect 11254 192574 11834 192658
rect 11254 192338 11426 192574
rect 11662 192338 11834 192574
rect 11254 156894 11834 192338
rect 11254 156658 11426 156894
rect 11662 156658 11834 156894
rect 11254 156574 11834 156658
rect 11254 156338 11426 156574
rect 11662 156338 11834 156574
rect 11254 120894 11834 156338
rect 11254 120658 11426 120894
rect 11662 120658 11834 120894
rect 11254 120574 11834 120658
rect 11254 120338 11426 120574
rect 11662 120338 11834 120574
rect 11254 84894 11834 120338
rect 11254 84658 11426 84894
rect 11662 84658 11834 84894
rect 11254 84574 11834 84658
rect 11254 84338 11426 84574
rect 11662 84338 11834 84574
rect 11254 48894 11834 84338
rect 11254 48658 11426 48894
rect 11662 48658 11834 48894
rect 11254 48574 11834 48658
rect 11254 48338 11426 48574
rect 11662 48338 11834 48574
rect 11254 12894 11834 48338
rect 11254 12658 11426 12894
rect 11662 12658 11834 12894
rect 11254 12574 11834 12658
rect 11254 12338 11426 12574
rect 11662 12338 11834 12574
rect -7506 -6102 -7334 -5866
rect -7098 -6102 -6926 -5866
rect -7506 -6186 -6926 -6102
rect -7506 -6422 -7334 -6186
rect -7098 -6422 -6926 -6186
rect -7506 -6434 -6926 -6422
rect 11254 -5866 11834 12338
rect 18814 705758 19394 705770
rect 18814 705522 18986 705758
rect 19222 705522 19394 705758
rect 18814 705438 19394 705522
rect 18814 705202 18986 705438
rect 19222 705202 19394 705438
rect 18814 668454 19394 705202
rect 18814 668218 18986 668454
rect 19222 668218 19394 668454
rect 18814 668134 19394 668218
rect 18814 667898 18986 668134
rect 19222 667898 19394 668134
rect 18814 632454 19394 667898
rect 18814 632218 18986 632454
rect 19222 632218 19394 632454
rect 18814 632134 19394 632218
rect 18814 631898 18986 632134
rect 19222 631898 19394 632134
rect 18814 596454 19394 631898
rect 18814 596218 18986 596454
rect 19222 596218 19394 596454
rect 18814 596134 19394 596218
rect 18814 595898 18986 596134
rect 19222 595898 19394 596134
rect 18814 560454 19394 595898
rect 18814 560218 18986 560454
rect 19222 560218 19394 560454
rect 18814 560134 19394 560218
rect 18814 559898 18986 560134
rect 19222 559898 19394 560134
rect 18814 524454 19394 559898
rect 18814 524218 18986 524454
rect 19222 524218 19394 524454
rect 18814 524134 19394 524218
rect 18814 523898 18986 524134
rect 19222 523898 19394 524134
rect 18814 488454 19394 523898
rect 18814 488218 18986 488454
rect 19222 488218 19394 488454
rect 18814 488134 19394 488218
rect 18814 487898 18986 488134
rect 19222 487898 19394 488134
rect 18814 452454 19394 487898
rect 18814 452218 18986 452454
rect 19222 452218 19394 452454
rect 18814 452134 19394 452218
rect 18814 451898 18986 452134
rect 19222 451898 19394 452134
rect 18814 416454 19394 451898
rect 18814 416218 18986 416454
rect 19222 416218 19394 416454
rect 18814 416134 19394 416218
rect 18814 415898 18986 416134
rect 19222 415898 19394 416134
rect 18814 380454 19394 415898
rect 18814 380218 18986 380454
rect 19222 380218 19394 380454
rect 18814 380134 19394 380218
rect 18814 379898 18986 380134
rect 19222 379898 19394 380134
rect 18814 344454 19394 379898
rect 18814 344218 18986 344454
rect 19222 344218 19394 344454
rect 18814 344134 19394 344218
rect 18814 343898 18986 344134
rect 19222 343898 19394 344134
rect 18814 308454 19394 343898
rect 18814 308218 18986 308454
rect 19222 308218 19394 308454
rect 18814 308134 19394 308218
rect 18814 307898 18986 308134
rect 19222 307898 19394 308134
rect 18814 272454 19394 307898
rect 18814 272218 18986 272454
rect 19222 272218 19394 272454
rect 18814 272134 19394 272218
rect 18814 271898 18986 272134
rect 19222 271898 19394 272134
rect 18814 236454 19394 271898
rect 18814 236218 18986 236454
rect 19222 236218 19394 236454
rect 18814 236134 19394 236218
rect 18814 235898 18986 236134
rect 19222 235898 19394 236134
rect 18814 200454 19394 235898
rect 18814 200218 18986 200454
rect 19222 200218 19394 200454
rect 18814 200134 19394 200218
rect 18814 199898 18986 200134
rect 19222 199898 19394 200134
rect 18814 164454 19394 199898
rect 18814 164218 18986 164454
rect 19222 164218 19394 164454
rect 18814 164134 19394 164218
rect 18814 163898 18986 164134
rect 19222 163898 19394 164134
rect 18814 128454 19394 163898
rect 18814 128218 18986 128454
rect 19222 128218 19394 128454
rect 18814 128134 19394 128218
rect 18814 127898 18986 128134
rect 19222 127898 19394 128134
rect 18814 92454 19394 127898
rect 18814 92218 18986 92454
rect 19222 92218 19394 92454
rect 18814 92134 19394 92218
rect 18814 91898 18986 92134
rect 19222 91898 19394 92134
rect 18814 56454 19394 91898
rect 18814 56218 18986 56454
rect 19222 56218 19394 56454
rect 18814 56134 19394 56218
rect 18814 55898 18986 56134
rect 19222 55898 19394 56134
rect 18814 20454 19394 55898
rect 18814 20218 18986 20454
rect 19222 20218 19394 20454
rect 18814 20134 19394 20218
rect 18814 19898 18986 20134
rect 19222 19898 19394 20134
rect 18814 -1266 19394 19898
rect 18814 -1502 18986 -1266
rect 19222 -1502 19394 -1266
rect 18814 -1586 19394 -1502
rect 18814 -1822 18986 -1586
rect 19222 -1822 19394 -1586
rect 18814 -1834 19394 -1822
rect 22294 671934 22874 707042
rect 22294 671698 22466 671934
rect 22702 671698 22874 671934
rect 22294 671614 22874 671698
rect 22294 671378 22466 671614
rect 22702 671378 22874 671614
rect 22294 635934 22874 671378
rect 22294 635698 22466 635934
rect 22702 635698 22874 635934
rect 22294 635614 22874 635698
rect 22294 635378 22466 635614
rect 22702 635378 22874 635614
rect 22294 599934 22874 635378
rect 22294 599698 22466 599934
rect 22702 599698 22874 599934
rect 22294 599614 22874 599698
rect 22294 599378 22466 599614
rect 22702 599378 22874 599614
rect 22294 563934 22874 599378
rect 22294 563698 22466 563934
rect 22702 563698 22874 563934
rect 22294 563614 22874 563698
rect 22294 563378 22466 563614
rect 22702 563378 22874 563614
rect 22294 527934 22874 563378
rect 22294 527698 22466 527934
rect 22702 527698 22874 527934
rect 22294 527614 22874 527698
rect 22294 527378 22466 527614
rect 22702 527378 22874 527614
rect 22294 491934 22874 527378
rect 22294 491698 22466 491934
rect 22702 491698 22874 491934
rect 22294 491614 22874 491698
rect 22294 491378 22466 491614
rect 22702 491378 22874 491614
rect 22294 455934 22874 491378
rect 22294 455698 22466 455934
rect 22702 455698 22874 455934
rect 22294 455614 22874 455698
rect 22294 455378 22466 455614
rect 22702 455378 22874 455614
rect 22294 419934 22874 455378
rect 22294 419698 22466 419934
rect 22702 419698 22874 419934
rect 22294 419614 22874 419698
rect 22294 419378 22466 419614
rect 22702 419378 22874 419614
rect 22294 383934 22874 419378
rect 22294 383698 22466 383934
rect 22702 383698 22874 383934
rect 22294 383614 22874 383698
rect 22294 383378 22466 383614
rect 22702 383378 22874 383614
rect 22294 347934 22874 383378
rect 22294 347698 22466 347934
rect 22702 347698 22874 347934
rect 22294 347614 22874 347698
rect 22294 347378 22466 347614
rect 22702 347378 22874 347614
rect 22294 311934 22874 347378
rect 22294 311698 22466 311934
rect 22702 311698 22874 311934
rect 22294 311614 22874 311698
rect 22294 311378 22466 311614
rect 22702 311378 22874 311614
rect 22294 275934 22874 311378
rect 22294 275698 22466 275934
rect 22702 275698 22874 275934
rect 22294 275614 22874 275698
rect 22294 275378 22466 275614
rect 22702 275378 22874 275614
rect 22294 239934 22874 275378
rect 22294 239698 22466 239934
rect 22702 239698 22874 239934
rect 22294 239614 22874 239698
rect 22294 239378 22466 239614
rect 22702 239378 22874 239614
rect 22294 203934 22874 239378
rect 22294 203698 22466 203934
rect 22702 203698 22874 203934
rect 22294 203614 22874 203698
rect 22294 203378 22466 203614
rect 22702 203378 22874 203614
rect 22294 167934 22874 203378
rect 22294 167698 22466 167934
rect 22702 167698 22874 167934
rect 22294 167614 22874 167698
rect 22294 167378 22466 167614
rect 22702 167378 22874 167614
rect 22294 131934 22874 167378
rect 22294 131698 22466 131934
rect 22702 131698 22874 131934
rect 22294 131614 22874 131698
rect 22294 131378 22466 131614
rect 22702 131378 22874 131614
rect 22294 95934 22874 131378
rect 22294 95698 22466 95934
rect 22702 95698 22874 95934
rect 22294 95614 22874 95698
rect 22294 95378 22466 95614
rect 22702 95378 22874 95614
rect 22294 59934 22874 95378
rect 22294 59698 22466 59934
rect 22702 59698 22874 59934
rect 22294 59614 22874 59698
rect 22294 59378 22466 59614
rect 22702 59378 22874 59614
rect 22294 23934 22874 59378
rect 22294 23698 22466 23934
rect 22702 23698 22874 23934
rect 22294 23614 22874 23698
rect 22294 23378 22466 23614
rect 22702 23378 22874 23614
rect 22294 -3106 22874 23378
rect 22294 -3342 22466 -3106
rect 22702 -3342 22874 -3106
rect 22294 -3426 22874 -3342
rect 22294 -3662 22466 -3426
rect 22702 -3662 22874 -3426
rect 22294 -3674 22874 -3662
rect 25774 675414 26354 708882
rect 25774 675178 25946 675414
rect 26182 675178 26354 675414
rect 25774 675094 26354 675178
rect 25774 674858 25946 675094
rect 26182 674858 26354 675094
rect 25774 639414 26354 674858
rect 25774 639178 25946 639414
rect 26182 639178 26354 639414
rect 25774 639094 26354 639178
rect 25774 638858 25946 639094
rect 26182 638858 26354 639094
rect 25774 603414 26354 638858
rect 25774 603178 25946 603414
rect 26182 603178 26354 603414
rect 25774 603094 26354 603178
rect 25774 602858 25946 603094
rect 26182 602858 26354 603094
rect 25774 567414 26354 602858
rect 25774 567178 25946 567414
rect 26182 567178 26354 567414
rect 25774 567094 26354 567178
rect 25774 566858 25946 567094
rect 26182 566858 26354 567094
rect 25774 531414 26354 566858
rect 25774 531178 25946 531414
rect 26182 531178 26354 531414
rect 25774 531094 26354 531178
rect 25774 530858 25946 531094
rect 26182 530858 26354 531094
rect 25774 495414 26354 530858
rect 25774 495178 25946 495414
rect 26182 495178 26354 495414
rect 25774 495094 26354 495178
rect 25774 494858 25946 495094
rect 26182 494858 26354 495094
rect 25774 459414 26354 494858
rect 25774 459178 25946 459414
rect 26182 459178 26354 459414
rect 25774 459094 26354 459178
rect 25774 458858 25946 459094
rect 26182 458858 26354 459094
rect 25774 423414 26354 458858
rect 25774 423178 25946 423414
rect 26182 423178 26354 423414
rect 25774 423094 26354 423178
rect 25774 422858 25946 423094
rect 26182 422858 26354 423094
rect 25774 387414 26354 422858
rect 25774 387178 25946 387414
rect 26182 387178 26354 387414
rect 25774 387094 26354 387178
rect 25774 386858 25946 387094
rect 26182 386858 26354 387094
rect 25774 351414 26354 386858
rect 25774 351178 25946 351414
rect 26182 351178 26354 351414
rect 25774 351094 26354 351178
rect 25774 350858 25946 351094
rect 26182 350858 26354 351094
rect 25774 315414 26354 350858
rect 25774 315178 25946 315414
rect 26182 315178 26354 315414
rect 25774 315094 26354 315178
rect 25774 314858 25946 315094
rect 26182 314858 26354 315094
rect 25774 279414 26354 314858
rect 25774 279178 25946 279414
rect 26182 279178 26354 279414
rect 25774 279094 26354 279178
rect 25774 278858 25946 279094
rect 26182 278858 26354 279094
rect 25774 243414 26354 278858
rect 25774 243178 25946 243414
rect 26182 243178 26354 243414
rect 25774 243094 26354 243178
rect 25774 242858 25946 243094
rect 26182 242858 26354 243094
rect 25774 207414 26354 242858
rect 25774 207178 25946 207414
rect 26182 207178 26354 207414
rect 25774 207094 26354 207178
rect 25774 206858 25946 207094
rect 26182 206858 26354 207094
rect 25774 171414 26354 206858
rect 25774 171178 25946 171414
rect 26182 171178 26354 171414
rect 25774 171094 26354 171178
rect 25774 170858 25946 171094
rect 26182 170858 26354 171094
rect 25774 135414 26354 170858
rect 25774 135178 25946 135414
rect 26182 135178 26354 135414
rect 25774 135094 26354 135178
rect 25774 134858 25946 135094
rect 26182 134858 26354 135094
rect 25774 99414 26354 134858
rect 25774 99178 25946 99414
rect 26182 99178 26354 99414
rect 25774 99094 26354 99178
rect 25774 98858 25946 99094
rect 26182 98858 26354 99094
rect 25774 63414 26354 98858
rect 25774 63178 25946 63414
rect 26182 63178 26354 63414
rect 25774 63094 26354 63178
rect 25774 62858 25946 63094
rect 26182 62858 26354 63094
rect 25774 27414 26354 62858
rect 25774 27178 25946 27414
rect 26182 27178 26354 27414
rect 25774 27094 26354 27178
rect 25774 26858 25946 27094
rect 26182 26858 26354 27094
rect 25774 -4946 26354 26858
rect 25774 -5182 25946 -4946
rect 26182 -5182 26354 -4946
rect 25774 -5266 26354 -5182
rect 25774 -5502 25946 -5266
rect 26182 -5502 26354 -5266
rect 25774 -5514 26354 -5502
rect 29254 678894 29834 710722
rect 47254 710358 47834 711290
rect 47254 710122 47426 710358
rect 47662 710122 47834 710358
rect 47254 710038 47834 710122
rect 47254 709802 47426 710038
rect 47662 709802 47834 710038
rect 43774 708518 44354 709450
rect 43774 708282 43946 708518
rect 44182 708282 44354 708518
rect 43774 708198 44354 708282
rect 43774 707962 43946 708198
rect 44182 707962 44354 708198
rect 40294 706678 40874 707610
rect 40294 706442 40466 706678
rect 40702 706442 40874 706678
rect 40294 706358 40874 706442
rect 40294 706122 40466 706358
rect 40702 706122 40874 706358
rect 29254 678658 29426 678894
rect 29662 678658 29834 678894
rect 29254 678574 29834 678658
rect 29254 678338 29426 678574
rect 29662 678338 29834 678574
rect 29254 642894 29834 678338
rect 29254 642658 29426 642894
rect 29662 642658 29834 642894
rect 29254 642574 29834 642658
rect 29254 642338 29426 642574
rect 29662 642338 29834 642574
rect 29254 606894 29834 642338
rect 29254 606658 29426 606894
rect 29662 606658 29834 606894
rect 29254 606574 29834 606658
rect 29254 606338 29426 606574
rect 29662 606338 29834 606574
rect 29254 570894 29834 606338
rect 29254 570658 29426 570894
rect 29662 570658 29834 570894
rect 29254 570574 29834 570658
rect 29254 570338 29426 570574
rect 29662 570338 29834 570574
rect 29254 534894 29834 570338
rect 29254 534658 29426 534894
rect 29662 534658 29834 534894
rect 29254 534574 29834 534658
rect 29254 534338 29426 534574
rect 29662 534338 29834 534574
rect 29254 498894 29834 534338
rect 29254 498658 29426 498894
rect 29662 498658 29834 498894
rect 29254 498574 29834 498658
rect 29254 498338 29426 498574
rect 29662 498338 29834 498574
rect 29254 462894 29834 498338
rect 29254 462658 29426 462894
rect 29662 462658 29834 462894
rect 29254 462574 29834 462658
rect 29254 462338 29426 462574
rect 29662 462338 29834 462574
rect 29254 426894 29834 462338
rect 29254 426658 29426 426894
rect 29662 426658 29834 426894
rect 29254 426574 29834 426658
rect 29254 426338 29426 426574
rect 29662 426338 29834 426574
rect 29254 390894 29834 426338
rect 29254 390658 29426 390894
rect 29662 390658 29834 390894
rect 29254 390574 29834 390658
rect 29254 390338 29426 390574
rect 29662 390338 29834 390574
rect 29254 354894 29834 390338
rect 29254 354658 29426 354894
rect 29662 354658 29834 354894
rect 29254 354574 29834 354658
rect 29254 354338 29426 354574
rect 29662 354338 29834 354574
rect 29254 318894 29834 354338
rect 29254 318658 29426 318894
rect 29662 318658 29834 318894
rect 29254 318574 29834 318658
rect 29254 318338 29426 318574
rect 29662 318338 29834 318574
rect 29254 282894 29834 318338
rect 29254 282658 29426 282894
rect 29662 282658 29834 282894
rect 29254 282574 29834 282658
rect 29254 282338 29426 282574
rect 29662 282338 29834 282574
rect 29254 246894 29834 282338
rect 29254 246658 29426 246894
rect 29662 246658 29834 246894
rect 29254 246574 29834 246658
rect 29254 246338 29426 246574
rect 29662 246338 29834 246574
rect 29254 210894 29834 246338
rect 29254 210658 29426 210894
rect 29662 210658 29834 210894
rect 29254 210574 29834 210658
rect 29254 210338 29426 210574
rect 29662 210338 29834 210574
rect 29254 174894 29834 210338
rect 29254 174658 29426 174894
rect 29662 174658 29834 174894
rect 29254 174574 29834 174658
rect 29254 174338 29426 174574
rect 29662 174338 29834 174574
rect 29254 138894 29834 174338
rect 29254 138658 29426 138894
rect 29662 138658 29834 138894
rect 29254 138574 29834 138658
rect 29254 138338 29426 138574
rect 29662 138338 29834 138574
rect 29254 102894 29834 138338
rect 29254 102658 29426 102894
rect 29662 102658 29834 102894
rect 29254 102574 29834 102658
rect 29254 102338 29426 102574
rect 29662 102338 29834 102574
rect 29254 66894 29834 102338
rect 29254 66658 29426 66894
rect 29662 66658 29834 66894
rect 29254 66574 29834 66658
rect 29254 66338 29426 66574
rect 29662 66338 29834 66574
rect 29254 30894 29834 66338
rect 29254 30658 29426 30894
rect 29662 30658 29834 30894
rect 29254 30574 29834 30658
rect 29254 30338 29426 30574
rect 29662 30338 29834 30574
rect 11254 -6102 11426 -5866
rect 11662 -6102 11834 -5866
rect 11254 -6186 11834 -6102
rect 11254 -6422 11426 -6186
rect 11662 -6422 11834 -6186
rect -8426 -7022 -8254 -6786
rect -8018 -7022 -7846 -6786
rect -8426 -7106 -7846 -7022
rect -8426 -7342 -8254 -7106
rect -8018 -7342 -7846 -7106
rect -8426 -7354 -7846 -7342
rect 11254 -7354 11834 -6422
rect 29254 -6786 29834 30338
rect 36814 704838 37394 705770
rect 36814 704602 36986 704838
rect 37222 704602 37394 704838
rect 36814 704518 37394 704602
rect 36814 704282 36986 704518
rect 37222 704282 37394 704518
rect 36814 686454 37394 704282
rect 36814 686218 36986 686454
rect 37222 686218 37394 686454
rect 36814 686134 37394 686218
rect 36814 685898 36986 686134
rect 37222 685898 37394 686134
rect 36814 650454 37394 685898
rect 36814 650218 36986 650454
rect 37222 650218 37394 650454
rect 36814 650134 37394 650218
rect 36814 649898 36986 650134
rect 37222 649898 37394 650134
rect 36814 614454 37394 649898
rect 36814 614218 36986 614454
rect 37222 614218 37394 614454
rect 36814 614134 37394 614218
rect 36814 613898 36986 614134
rect 37222 613898 37394 614134
rect 36814 578454 37394 613898
rect 36814 578218 36986 578454
rect 37222 578218 37394 578454
rect 36814 578134 37394 578218
rect 36814 577898 36986 578134
rect 37222 577898 37394 578134
rect 36814 542454 37394 577898
rect 36814 542218 36986 542454
rect 37222 542218 37394 542454
rect 36814 542134 37394 542218
rect 36814 541898 36986 542134
rect 37222 541898 37394 542134
rect 36814 506454 37394 541898
rect 36814 506218 36986 506454
rect 37222 506218 37394 506454
rect 36814 506134 37394 506218
rect 36814 505898 36986 506134
rect 37222 505898 37394 506134
rect 36814 470454 37394 505898
rect 36814 470218 36986 470454
rect 37222 470218 37394 470454
rect 36814 470134 37394 470218
rect 36814 469898 36986 470134
rect 37222 469898 37394 470134
rect 36814 434454 37394 469898
rect 36814 434218 36986 434454
rect 37222 434218 37394 434454
rect 36814 434134 37394 434218
rect 36814 433898 36986 434134
rect 37222 433898 37394 434134
rect 36814 398454 37394 433898
rect 36814 398218 36986 398454
rect 37222 398218 37394 398454
rect 36814 398134 37394 398218
rect 36814 397898 36986 398134
rect 37222 397898 37394 398134
rect 36814 362454 37394 397898
rect 36814 362218 36986 362454
rect 37222 362218 37394 362454
rect 36814 362134 37394 362218
rect 36814 361898 36986 362134
rect 37222 361898 37394 362134
rect 36814 326454 37394 361898
rect 36814 326218 36986 326454
rect 37222 326218 37394 326454
rect 36814 326134 37394 326218
rect 36814 325898 36986 326134
rect 37222 325898 37394 326134
rect 36814 290454 37394 325898
rect 36814 290218 36986 290454
rect 37222 290218 37394 290454
rect 36814 290134 37394 290218
rect 36814 289898 36986 290134
rect 37222 289898 37394 290134
rect 36814 254454 37394 289898
rect 36814 254218 36986 254454
rect 37222 254218 37394 254454
rect 36814 254134 37394 254218
rect 36814 253898 36986 254134
rect 37222 253898 37394 254134
rect 36814 218454 37394 253898
rect 36814 218218 36986 218454
rect 37222 218218 37394 218454
rect 36814 218134 37394 218218
rect 36814 217898 36986 218134
rect 37222 217898 37394 218134
rect 36814 182454 37394 217898
rect 36814 182218 36986 182454
rect 37222 182218 37394 182454
rect 36814 182134 37394 182218
rect 36814 181898 36986 182134
rect 37222 181898 37394 182134
rect 36814 146454 37394 181898
rect 36814 146218 36986 146454
rect 37222 146218 37394 146454
rect 36814 146134 37394 146218
rect 36814 145898 36986 146134
rect 37222 145898 37394 146134
rect 36814 110454 37394 145898
rect 36814 110218 36986 110454
rect 37222 110218 37394 110454
rect 36814 110134 37394 110218
rect 36814 109898 36986 110134
rect 37222 109898 37394 110134
rect 36814 74454 37394 109898
rect 36814 74218 36986 74454
rect 37222 74218 37394 74454
rect 36814 74134 37394 74218
rect 36814 73898 36986 74134
rect 37222 73898 37394 74134
rect 36814 38454 37394 73898
rect 36814 38218 36986 38454
rect 37222 38218 37394 38454
rect 36814 38134 37394 38218
rect 36814 37898 36986 38134
rect 37222 37898 37394 38134
rect 36814 2454 37394 37898
rect 36814 2218 36986 2454
rect 37222 2218 37394 2454
rect 36814 2134 37394 2218
rect 36814 1898 36986 2134
rect 37222 1898 37394 2134
rect 36814 -346 37394 1898
rect 36814 -582 36986 -346
rect 37222 -582 37394 -346
rect 36814 -666 37394 -582
rect 36814 -902 36986 -666
rect 37222 -902 37394 -666
rect 36814 -1834 37394 -902
rect 40294 689934 40874 706122
rect 40294 689698 40466 689934
rect 40702 689698 40874 689934
rect 40294 689614 40874 689698
rect 40294 689378 40466 689614
rect 40702 689378 40874 689614
rect 40294 653934 40874 689378
rect 40294 653698 40466 653934
rect 40702 653698 40874 653934
rect 40294 653614 40874 653698
rect 40294 653378 40466 653614
rect 40702 653378 40874 653614
rect 40294 617934 40874 653378
rect 40294 617698 40466 617934
rect 40702 617698 40874 617934
rect 40294 617614 40874 617698
rect 40294 617378 40466 617614
rect 40702 617378 40874 617614
rect 40294 581934 40874 617378
rect 40294 581698 40466 581934
rect 40702 581698 40874 581934
rect 40294 581614 40874 581698
rect 40294 581378 40466 581614
rect 40702 581378 40874 581614
rect 40294 545934 40874 581378
rect 40294 545698 40466 545934
rect 40702 545698 40874 545934
rect 40294 545614 40874 545698
rect 40294 545378 40466 545614
rect 40702 545378 40874 545614
rect 40294 509934 40874 545378
rect 40294 509698 40466 509934
rect 40702 509698 40874 509934
rect 40294 509614 40874 509698
rect 40294 509378 40466 509614
rect 40702 509378 40874 509614
rect 40294 473934 40874 509378
rect 40294 473698 40466 473934
rect 40702 473698 40874 473934
rect 40294 473614 40874 473698
rect 40294 473378 40466 473614
rect 40702 473378 40874 473614
rect 40294 437934 40874 473378
rect 40294 437698 40466 437934
rect 40702 437698 40874 437934
rect 40294 437614 40874 437698
rect 40294 437378 40466 437614
rect 40702 437378 40874 437614
rect 40294 401934 40874 437378
rect 40294 401698 40466 401934
rect 40702 401698 40874 401934
rect 40294 401614 40874 401698
rect 40294 401378 40466 401614
rect 40702 401378 40874 401614
rect 40294 365934 40874 401378
rect 40294 365698 40466 365934
rect 40702 365698 40874 365934
rect 40294 365614 40874 365698
rect 40294 365378 40466 365614
rect 40702 365378 40874 365614
rect 40294 329934 40874 365378
rect 40294 329698 40466 329934
rect 40702 329698 40874 329934
rect 40294 329614 40874 329698
rect 40294 329378 40466 329614
rect 40702 329378 40874 329614
rect 40294 293934 40874 329378
rect 40294 293698 40466 293934
rect 40702 293698 40874 293934
rect 40294 293614 40874 293698
rect 40294 293378 40466 293614
rect 40702 293378 40874 293614
rect 40294 257934 40874 293378
rect 40294 257698 40466 257934
rect 40702 257698 40874 257934
rect 40294 257614 40874 257698
rect 40294 257378 40466 257614
rect 40702 257378 40874 257614
rect 40294 221934 40874 257378
rect 40294 221698 40466 221934
rect 40702 221698 40874 221934
rect 40294 221614 40874 221698
rect 40294 221378 40466 221614
rect 40702 221378 40874 221614
rect 40294 185934 40874 221378
rect 40294 185698 40466 185934
rect 40702 185698 40874 185934
rect 40294 185614 40874 185698
rect 40294 185378 40466 185614
rect 40702 185378 40874 185614
rect 40294 149934 40874 185378
rect 40294 149698 40466 149934
rect 40702 149698 40874 149934
rect 40294 149614 40874 149698
rect 40294 149378 40466 149614
rect 40702 149378 40874 149614
rect 40294 113934 40874 149378
rect 40294 113698 40466 113934
rect 40702 113698 40874 113934
rect 40294 113614 40874 113698
rect 40294 113378 40466 113614
rect 40702 113378 40874 113614
rect 40294 77934 40874 113378
rect 40294 77698 40466 77934
rect 40702 77698 40874 77934
rect 40294 77614 40874 77698
rect 40294 77378 40466 77614
rect 40702 77378 40874 77614
rect 40294 41934 40874 77378
rect 40294 41698 40466 41934
rect 40702 41698 40874 41934
rect 40294 41614 40874 41698
rect 40294 41378 40466 41614
rect 40702 41378 40874 41614
rect 40294 5934 40874 41378
rect 40294 5698 40466 5934
rect 40702 5698 40874 5934
rect 40294 5614 40874 5698
rect 40294 5378 40466 5614
rect 40702 5378 40874 5614
rect 40294 -2186 40874 5378
rect 40294 -2422 40466 -2186
rect 40702 -2422 40874 -2186
rect 40294 -2506 40874 -2422
rect 40294 -2742 40466 -2506
rect 40702 -2742 40874 -2506
rect 40294 -3674 40874 -2742
rect 43774 693414 44354 707962
rect 43774 693178 43946 693414
rect 44182 693178 44354 693414
rect 43774 693094 44354 693178
rect 43774 692858 43946 693094
rect 44182 692858 44354 693094
rect 43774 657414 44354 692858
rect 43774 657178 43946 657414
rect 44182 657178 44354 657414
rect 43774 657094 44354 657178
rect 43774 656858 43946 657094
rect 44182 656858 44354 657094
rect 43774 621414 44354 656858
rect 43774 621178 43946 621414
rect 44182 621178 44354 621414
rect 43774 621094 44354 621178
rect 43774 620858 43946 621094
rect 44182 620858 44354 621094
rect 43774 585414 44354 620858
rect 43774 585178 43946 585414
rect 44182 585178 44354 585414
rect 43774 585094 44354 585178
rect 43774 584858 43946 585094
rect 44182 584858 44354 585094
rect 43774 549414 44354 584858
rect 43774 549178 43946 549414
rect 44182 549178 44354 549414
rect 43774 549094 44354 549178
rect 43774 548858 43946 549094
rect 44182 548858 44354 549094
rect 43774 513414 44354 548858
rect 43774 513178 43946 513414
rect 44182 513178 44354 513414
rect 43774 513094 44354 513178
rect 43774 512858 43946 513094
rect 44182 512858 44354 513094
rect 43774 477414 44354 512858
rect 43774 477178 43946 477414
rect 44182 477178 44354 477414
rect 43774 477094 44354 477178
rect 43774 476858 43946 477094
rect 44182 476858 44354 477094
rect 43774 441414 44354 476858
rect 43774 441178 43946 441414
rect 44182 441178 44354 441414
rect 43774 441094 44354 441178
rect 43774 440858 43946 441094
rect 44182 440858 44354 441094
rect 43774 405414 44354 440858
rect 43774 405178 43946 405414
rect 44182 405178 44354 405414
rect 43774 405094 44354 405178
rect 43774 404858 43946 405094
rect 44182 404858 44354 405094
rect 43774 369414 44354 404858
rect 43774 369178 43946 369414
rect 44182 369178 44354 369414
rect 43774 369094 44354 369178
rect 43774 368858 43946 369094
rect 44182 368858 44354 369094
rect 43774 333414 44354 368858
rect 43774 333178 43946 333414
rect 44182 333178 44354 333414
rect 43774 333094 44354 333178
rect 43774 332858 43946 333094
rect 44182 332858 44354 333094
rect 43774 297414 44354 332858
rect 43774 297178 43946 297414
rect 44182 297178 44354 297414
rect 43774 297094 44354 297178
rect 43774 296858 43946 297094
rect 44182 296858 44354 297094
rect 43774 261414 44354 296858
rect 43774 261178 43946 261414
rect 44182 261178 44354 261414
rect 43774 261094 44354 261178
rect 43774 260858 43946 261094
rect 44182 260858 44354 261094
rect 43774 225414 44354 260858
rect 43774 225178 43946 225414
rect 44182 225178 44354 225414
rect 43774 225094 44354 225178
rect 43774 224858 43946 225094
rect 44182 224858 44354 225094
rect 43774 189414 44354 224858
rect 43774 189178 43946 189414
rect 44182 189178 44354 189414
rect 43774 189094 44354 189178
rect 43774 188858 43946 189094
rect 44182 188858 44354 189094
rect 43774 153414 44354 188858
rect 43774 153178 43946 153414
rect 44182 153178 44354 153414
rect 43774 153094 44354 153178
rect 43774 152858 43946 153094
rect 44182 152858 44354 153094
rect 43774 117414 44354 152858
rect 43774 117178 43946 117414
rect 44182 117178 44354 117414
rect 43774 117094 44354 117178
rect 43774 116858 43946 117094
rect 44182 116858 44354 117094
rect 43774 81414 44354 116858
rect 43774 81178 43946 81414
rect 44182 81178 44354 81414
rect 43774 81094 44354 81178
rect 43774 80858 43946 81094
rect 44182 80858 44354 81094
rect 43774 45414 44354 80858
rect 43774 45178 43946 45414
rect 44182 45178 44354 45414
rect 43774 45094 44354 45178
rect 43774 44858 43946 45094
rect 44182 44858 44354 45094
rect 43774 9414 44354 44858
rect 43774 9178 43946 9414
rect 44182 9178 44354 9414
rect 43774 9094 44354 9178
rect 43774 8858 43946 9094
rect 44182 8858 44354 9094
rect 43774 -4026 44354 8858
rect 43774 -4262 43946 -4026
rect 44182 -4262 44354 -4026
rect 43774 -4346 44354 -4262
rect 43774 -4582 43946 -4346
rect 44182 -4582 44354 -4346
rect 43774 -5514 44354 -4582
rect 47254 696894 47834 709802
rect 65254 711278 65834 711290
rect 65254 711042 65426 711278
rect 65662 711042 65834 711278
rect 65254 710958 65834 711042
rect 65254 710722 65426 710958
rect 65662 710722 65834 710958
rect 61774 709438 62354 709450
rect 61774 709202 61946 709438
rect 62182 709202 62354 709438
rect 61774 709118 62354 709202
rect 61774 708882 61946 709118
rect 62182 708882 62354 709118
rect 58294 707598 58874 707610
rect 58294 707362 58466 707598
rect 58702 707362 58874 707598
rect 58294 707278 58874 707362
rect 58294 707042 58466 707278
rect 58702 707042 58874 707278
rect 47254 696658 47426 696894
rect 47662 696658 47834 696894
rect 47254 696574 47834 696658
rect 47254 696338 47426 696574
rect 47662 696338 47834 696574
rect 47254 660894 47834 696338
rect 47254 660658 47426 660894
rect 47662 660658 47834 660894
rect 47254 660574 47834 660658
rect 47254 660338 47426 660574
rect 47662 660338 47834 660574
rect 47254 624894 47834 660338
rect 47254 624658 47426 624894
rect 47662 624658 47834 624894
rect 47254 624574 47834 624658
rect 47254 624338 47426 624574
rect 47662 624338 47834 624574
rect 47254 588894 47834 624338
rect 47254 588658 47426 588894
rect 47662 588658 47834 588894
rect 47254 588574 47834 588658
rect 47254 588338 47426 588574
rect 47662 588338 47834 588574
rect 47254 552894 47834 588338
rect 47254 552658 47426 552894
rect 47662 552658 47834 552894
rect 47254 552574 47834 552658
rect 47254 552338 47426 552574
rect 47662 552338 47834 552574
rect 47254 516894 47834 552338
rect 47254 516658 47426 516894
rect 47662 516658 47834 516894
rect 47254 516574 47834 516658
rect 47254 516338 47426 516574
rect 47662 516338 47834 516574
rect 47254 480894 47834 516338
rect 47254 480658 47426 480894
rect 47662 480658 47834 480894
rect 47254 480574 47834 480658
rect 47254 480338 47426 480574
rect 47662 480338 47834 480574
rect 47254 444894 47834 480338
rect 47254 444658 47426 444894
rect 47662 444658 47834 444894
rect 47254 444574 47834 444658
rect 47254 444338 47426 444574
rect 47662 444338 47834 444574
rect 47254 408894 47834 444338
rect 47254 408658 47426 408894
rect 47662 408658 47834 408894
rect 47254 408574 47834 408658
rect 47254 408338 47426 408574
rect 47662 408338 47834 408574
rect 47254 372894 47834 408338
rect 47254 372658 47426 372894
rect 47662 372658 47834 372894
rect 47254 372574 47834 372658
rect 47254 372338 47426 372574
rect 47662 372338 47834 372574
rect 47254 336894 47834 372338
rect 47254 336658 47426 336894
rect 47662 336658 47834 336894
rect 47254 336574 47834 336658
rect 47254 336338 47426 336574
rect 47662 336338 47834 336574
rect 47254 300894 47834 336338
rect 47254 300658 47426 300894
rect 47662 300658 47834 300894
rect 47254 300574 47834 300658
rect 47254 300338 47426 300574
rect 47662 300338 47834 300574
rect 47254 264894 47834 300338
rect 47254 264658 47426 264894
rect 47662 264658 47834 264894
rect 47254 264574 47834 264658
rect 47254 264338 47426 264574
rect 47662 264338 47834 264574
rect 47254 228894 47834 264338
rect 47254 228658 47426 228894
rect 47662 228658 47834 228894
rect 47254 228574 47834 228658
rect 47254 228338 47426 228574
rect 47662 228338 47834 228574
rect 47254 192894 47834 228338
rect 47254 192658 47426 192894
rect 47662 192658 47834 192894
rect 47254 192574 47834 192658
rect 47254 192338 47426 192574
rect 47662 192338 47834 192574
rect 47254 156894 47834 192338
rect 47254 156658 47426 156894
rect 47662 156658 47834 156894
rect 47254 156574 47834 156658
rect 47254 156338 47426 156574
rect 47662 156338 47834 156574
rect 47254 120894 47834 156338
rect 47254 120658 47426 120894
rect 47662 120658 47834 120894
rect 47254 120574 47834 120658
rect 47254 120338 47426 120574
rect 47662 120338 47834 120574
rect 47254 84894 47834 120338
rect 47254 84658 47426 84894
rect 47662 84658 47834 84894
rect 47254 84574 47834 84658
rect 47254 84338 47426 84574
rect 47662 84338 47834 84574
rect 47254 48894 47834 84338
rect 47254 48658 47426 48894
rect 47662 48658 47834 48894
rect 47254 48574 47834 48658
rect 47254 48338 47426 48574
rect 47662 48338 47834 48574
rect 47254 12894 47834 48338
rect 47254 12658 47426 12894
rect 47662 12658 47834 12894
rect 47254 12574 47834 12658
rect 47254 12338 47426 12574
rect 47662 12338 47834 12574
rect 29254 -7022 29426 -6786
rect 29662 -7022 29834 -6786
rect 29254 -7106 29834 -7022
rect 29254 -7342 29426 -7106
rect 29662 -7342 29834 -7106
rect 29254 -7354 29834 -7342
rect 47254 -5866 47834 12338
rect 54814 705758 55394 705770
rect 54814 705522 54986 705758
rect 55222 705522 55394 705758
rect 54814 705438 55394 705522
rect 54814 705202 54986 705438
rect 55222 705202 55394 705438
rect 54814 668454 55394 705202
rect 54814 668218 54986 668454
rect 55222 668218 55394 668454
rect 54814 668134 55394 668218
rect 54814 667898 54986 668134
rect 55222 667898 55394 668134
rect 54814 632454 55394 667898
rect 54814 632218 54986 632454
rect 55222 632218 55394 632454
rect 54814 632134 55394 632218
rect 54814 631898 54986 632134
rect 55222 631898 55394 632134
rect 54814 596454 55394 631898
rect 54814 596218 54986 596454
rect 55222 596218 55394 596454
rect 54814 596134 55394 596218
rect 54814 595898 54986 596134
rect 55222 595898 55394 596134
rect 54814 560454 55394 595898
rect 54814 560218 54986 560454
rect 55222 560218 55394 560454
rect 54814 560134 55394 560218
rect 54814 559898 54986 560134
rect 55222 559898 55394 560134
rect 54814 524454 55394 559898
rect 54814 524218 54986 524454
rect 55222 524218 55394 524454
rect 54814 524134 55394 524218
rect 54814 523898 54986 524134
rect 55222 523898 55394 524134
rect 54814 488454 55394 523898
rect 54814 488218 54986 488454
rect 55222 488218 55394 488454
rect 54814 488134 55394 488218
rect 54814 487898 54986 488134
rect 55222 487898 55394 488134
rect 54814 452454 55394 487898
rect 54814 452218 54986 452454
rect 55222 452218 55394 452454
rect 54814 452134 55394 452218
rect 54814 451898 54986 452134
rect 55222 451898 55394 452134
rect 54814 416454 55394 451898
rect 54814 416218 54986 416454
rect 55222 416218 55394 416454
rect 54814 416134 55394 416218
rect 54814 415898 54986 416134
rect 55222 415898 55394 416134
rect 54814 380454 55394 415898
rect 54814 380218 54986 380454
rect 55222 380218 55394 380454
rect 54814 380134 55394 380218
rect 54814 379898 54986 380134
rect 55222 379898 55394 380134
rect 54814 344454 55394 379898
rect 54814 344218 54986 344454
rect 55222 344218 55394 344454
rect 54814 344134 55394 344218
rect 54814 343898 54986 344134
rect 55222 343898 55394 344134
rect 54814 308454 55394 343898
rect 54814 308218 54986 308454
rect 55222 308218 55394 308454
rect 54814 308134 55394 308218
rect 54814 307898 54986 308134
rect 55222 307898 55394 308134
rect 54814 272454 55394 307898
rect 54814 272218 54986 272454
rect 55222 272218 55394 272454
rect 54814 272134 55394 272218
rect 54814 271898 54986 272134
rect 55222 271898 55394 272134
rect 54814 236454 55394 271898
rect 54814 236218 54986 236454
rect 55222 236218 55394 236454
rect 54814 236134 55394 236218
rect 54814 235898 54986 236134
rect 55222 235898 55394 236134
rect 54814 200454 55394 235898
rect 54814 200218 54986 200454
rect 55222 200218 55394 200454
rect 54814 200134 55394 200218
rect 54814 199898 54986 200134
rect 55222 199898 55394 200134
rect 54814 164454 55394 199898
rect 54814 164218 54986 164454
rect 55222 164218 55394 164454
rect 54814 164134 55394 164218
rect 54814 163898 54986 164134
rect 55222 163898 55394 164134
rect 54814 128454 55394 163898
rect 54814 128218 54986 128454
rect 55222 128218 55394 128454
rect 54814 128134 55394 128218
rect 54814 127898 54986 128134
rect 55222 127898 55394 128134
rect 54814 92454 55394 127898
rect 54814 92218 54986 92454
rect 55222 92218 55394 92454
rect 54814 92134 55394 92218
rect 54814 91898 54986 92134
rect 55222 91898 55394 92134
rect 54814 56454 55394 91898
rect 54814 56218 54986 56454
rect 55222 56218 55394 56454
rect 54814 56134 55394 56218
rect 54814 55898 54986 56134
rect 55222 55898 55394 56134
rect 54814 20454 55394 55898
rect 54814 20218 54986 20454
rect 55222 20218 55394 20454
rect 54814 20134 55394 20218
rect 54814 19898 54986 20134
rect 55222 19898 55394 20134
rect 54814 -1266 55394 19898
rect 54814 -1502 54986 -1266
rect 55222 -1502 55394 -1266
rect 54814 -1586 55394 -1502
rect 54814 -1822 54986 -1586
rect 55222 -1822 55394 -1586
rect 54814 -1834 55394 -1822
rect 58294 671934 58874 707042
rect 58294 671698 58466 671934
rect 58702 671698 58874 671934
rect 58294 671614 58874 671698
rect 58294 671378 58466 671614
rect 58702 671378 58874 671614
rect 58294 635934 58874 671378
rect 58294 635698 58466 635934
rect 58702 635698 58874 635934
rect 58294 635614 58874 635698
rect 58294 635378 58466 635614
rect 58702 635378 58874 635614
rect 58294 599934 58874 635378
rect 58294 599698 58466 599934
rect 58702 599698 58874 599934
rect 58294 599614 58874 599698
rect 58294 599378 58466 599614
rect 58702 599378 58874 599614
rect 58294 563934 58874 599378
rect 58294 563698 58466 563934
rect 58702 563698 58874 563934
rect 58294 563614 58874 563698
rect 58294 563378 58466 563614
rect 58702 563378 58874 563614
rect 58294 527934 58874 563378
rect 58294 527698 58466 527934
rect 58702 527698 58874 527934
rect 58294 527614 58874 527698
rect 58294 527378 58466 527614
rect 58702 527378 58874 527614
rect 58294 491934 58874 527378
rect 58294 491698 58466 491934
rect 58702 491698 58874 491934
rect 58294 491614 58874 491698
rect 58294 491378 58466 491614
rect 58702 491378 58874 491614
rect 58294 455934 58874 491378
rect 58294 455698 58466 455934
rect 58702 455698 58874 455934
rect 58294 455614 58874 455698
rect 58294 455378 58466 455614
rect 58702 455378 58874 455614
rect 58294 419934 58874 455378
rect 58294 419698 58466 419934
rect 58702 419698 58874 419934
rect 58294 419614 58874 419698
rect 58294 419378 58466 419614
rect 58702 419378 58874 419614
rect 58294 383934 58874 419378
rect 58294 383698 58466 383934
rect 58702 383698 58874 383934
rect 58294 383614 58874 383698
rect 58294 383378 58466 383614
rect 58702 383378 58874 383614
rect 58294 347934 58874 383378
rect 58294 347698 58466 347934
rect 58702 347698 58874 347934
rect 58294 347614 58874 347698
rect 58294 347378 58466 347614
rect 58702 347378 58874 347614
rect 58294 311934 58874 347378
rect 58294 311698 58466 311934
rect 58702 311698 58874 311934
rect 58294 311614 58874 311698
rect 58294 311378 58466 311614
rect 58702 311378 58874 311614
rect 58294 275934 58874 311378
rect 58294 275698 58466 275934
rect 58702 275698 58874 275934
rect 58294 275614 58874 275698
rect 58294 275378 58466 275614
rect 58702 275378 58874 275614
rect 58294 239934 58874 275378
rect 58294 239698 58466 239934
rect 58702 239698 58874 239934
rect 58294 239614 58874 239698
rect 58294 239378 58466 239614
rect 58702 239378 58874 239614
rect 58294 203934 58874 239378
rect 58294 203698 58466 203934
rect 58702 203698 58874 203934
rect 58294 203614 58874 203698
rect 58294 203378 58466 203614
rect 58702 203378 58874 203614
rect 58294 167934 58874 203378
rect 58294 167698 58466 167934
rect 58702 167698 58874 167934
rect 58294 167614 58874 167698
rect 58294 167378 58466 167614
rect 58702 167378 58874 167614
rect 58294 131934 58874 167378
rect 58294 131698 58466 131934
rect 58702 131698 58874 131934
rect 58294 131614 58874 131698
rect 58294 131378 58466 131614
rect 58702 131378 58874 131614
rect 58294 95934 58874 131378
rect 58294 95698 58466 95934
rect 58702 95698 58874 95934
rect 58294 95614 58874 95698
rect 58294 95378 58466 95614
rect 58702 95378 58874 95614
rect 58294 59934 58874 95378
rect 58294 59698 58466 59934
rect 58702 59698 58874 59934
rect 58294 59614 58874 59698
rect 58294 59378 58466 59614
rect 58702 59378 58874 59614
rect 58294 23934 58874 59378
rect 58294 23698 58466 23934
rect 58702 23698 58874 23934
rect 58294 23614 58874 23698
rect 58294 23378 58466 23614
rect 58702 23378 58874 23614
rect 58294 -3106 58874 23378
rect 58294 -3342 58466 -3106
rect 58702 -3342 58874 -3106
rect 58294 -3426 58874 -3342
rect 58294 -3662 58466 -3426
rect 58702 -3662 58874 -3426
rect 58294 -3674 58874 -3662
rect 61774 675414 62354 708882
rect 61774 675178 61946 675414
rect 62182 675178 62354 675414
rect 61774 675094 62354 675178
rect 61774 674858 61946 675094
rect 62182 674858 62354 675094
rect 61774 639414 62354 674858
rect 61774 639178 61946 639414
rect 62182 639178 62354 639414
rect 61774 639094 62354 639178
rect 61774 638858 61946 639094
rect 62182 638858 62354 639094
rect 61774 603414 62354 638858
rect 61774 603178 61946 603414
rect 62182 603178 62354 603414
rect 61774 603094 62354 603178
rect 61774 602858 61946 603094
rect 62182 602858 62354 603094
rect 61774 567414 62354 602858
rect 61774 567178 61946 567414
rect 62182 567178 62354 567414
rect 61774 567094 62354 567178
rect 61774 566858 61946 567094
rect 62182 566858 62354 567094
rect 61774 531414 62354 566858
rect 61774 531178 61946 531414
rect 62182 531178 62354 531414
rect 61774 531094 62354 531178
rect 61774 530858 61946 531094
rect 62182 530858 62354 531094
rect 61774 495414 62354 530858
rect 61774 495178 61946 495414
rect 62182 495178 62354 495414
rect 61774 495094 62354 495178
rect 61774 494858 61946 495094
rect 62182 494858 62354 495094
rect 61774 459414 62354 494858
rect 61774 459178 61946 459414
rect 62182 459178 62354 459414
rect 61774 459094 62354 459178
rect 61774 458858 61946 459094
rect 62182 458858 62354 459094
rect 61774 423414 62354 458858
rect 61774 423178 61946 423414
rect 62182 423178 62354 423414
rect 61774 423094 62354 423178
rect 61774 422858 61946 423094
rect 62182 422858 62354 423094
rect 61774 387414 62354 422858
rect 61774 387178 61946 387414
rect 62182 387178 62354 387414
rect 61774 387094 62354 387178
rect 61774 386858 61946 387094
rect 62182 386858 62354 387094
rect 61774 351414 62354 386858
rect 61774 351178 61946 351414
rect 62182 351178 62354 351414
rect 61774 351094 62354 351178
rect 61774 350858 61946 351094
rect 62182 350858 62354 351094
rect 61774 315414 62354 350858
rect 61774 315178 61946 315414
rect 62182 315178 62354 315414
rect 61774 315094 62354 315178
rect 61774 314858 61946 315094
rect 62182 314858 62354 315094
rect 61774 279414 62354 314858
rect 61774 279178 61946 279414
rect 62182 279178 62354 279414
rect 61774 279094 62354 279178
rect 61774 278858 61946 279094
rect 62182 278858 62354 279094
rect 61774 243414 62354 278858
rect 61774 243178 61946 243414
rect 62182 243178 62354 243414
rect 61774 243094 62354 243178
rect 61774 242858 61946 243094
rect 62182 242858 62354 243094
rect 61774 207414 62354 242858
rect 61774 207178 61946 207414
rect 62182 207178 62354 207414
rect 61774 207094 62354 207178
rect 61774 206858 61946 207094
rect 62182 206858 62354 207094
rect 61774 171414 62354 206858
rect 61774 171178 61946 171414
rect 62182 171178 62354 171414
rect 61774 171094 62354 171178
rect 61774 170858 61946 171094
rect 62182 170858 62354 171094
rect 61774 135414 62354 170858
rect 61774 135178 61946 135414
rect 62182 135178 62354 135414
rect 61774 135094 62354 135178
rect 61774 134858 61946 135094
rect 62182 134858 62354 135094
rect 61774 99414 62354 134858
rect 61774 99178 61946 99414
rect 62182 99178 62354 99414
rect 61774 99094 62354 99178
rect 61774 98858 61946 99094
rect 62182 98858 62354 99094
rect 61774 63414 62354 98858
rect 61774 63178 61946 63414
rect 62182 63178 62354 63414
rect 61774 63094 62354 63178
rect 61774 62858 61946 63094
rect 62182 62858 62354 63094
rect 61774 27414 62354 62858
rect 61774 27178 61946 27414
rect 62182 27178 62354 27414
rect 61774 27094 62354 27178
rect 61774 26858 61946 27094
rect 62182 26858 62354 27094
rect 61774 -4946 62354 26858
rect 61774 -5182 61946 -4946
rect 62182 -5182 62354 -4946
rect 61774 -5266 62354 -5182
rect 61774 -5502 61946 -5266
rect 62182 -5502 62354 -5266
rect 61774 -5514 62354 -5502
rect 65254 678894 65834 710722
rect 83254 710358 83834 711290
rect 83254 710122 83426 710358
rect 83662 710122 83834 710358
rect 83254 710038 83834 710122
rect 83254 709802 83426 710038
rect 83662 709802 83834 710038
rect 79774 708518 80354 709450
rect 79774 708282 79946 708518
rect 80182 708282 80354 708518
rect 79774 708198 80354 708282
rect 79774 707962 79946 708198
rect 80182 707962 80354 708198
rect 76294 706678 76874 707610
rect 76294 706442 76466 706678
rect 76702 706442 76874 706678
rect 76294 706358 76874 706442
rect 76294 706122 76466 706358
rect 76702 706122 76874 706358
rect 65254 678658 65426 678894
rect 65662 678658 65834 678894
rect 65254 678574 65834 678658
rect 65254 678338 65426 678574
rect 65662 678338 65834 678574
rect 65254 642894 65834 678338
rect 65254 642658 65426 642894
rect 65662 642658 65834 642894
rect 65254 642574 65834 642658
rect 65254 642338 65426 642574
rect 65662 642338 65834 642574
rect 65254 606894 65834 642338
rect 65254 606658 65426 606894
rect 65662 606658 65834 606894
rect 65254 606574 65834 606658
rect 65254 606338 65426 606574
rect 65662 606338 65834 606574
rect 65254 570894 65834 606338
rect 65254 570658 65426 570894
rect 65662 570658 65834 570894
rect 65254 570574 65834 570658
rect 65254 570338 65426 570574
rect 65662 570338 65834 570574
rect 65254 534894 65834 570338
rect 65254 534658 65426 534894
rect 65662 534658 65834 534894
rect 65254 534574 65834 534658
rect 65254 534338 65426 534574
rect 65662 534338 65834 534574
rect 65254 498894 65834 534338
rect 65254 498658 65426 498894
rect 65662 498658 65834 498894
rect 65254 498574 65834 498658
rect 65254 498338 65426 498574
rect 65662 498338 65834 498574
rect 65254 462894 65834 498338
rect 65254 462658 65426 462894
rect 65662 462658 65834 462894
rect 65254 462574 65834 462658
rect 65254 462338 65426 462574
rect 65662 462338 65834 462574
rect 65254 426894 65834 462338
rect 65254 426658 65426 426894
rect 65662 426658 65834 426894
rect 65254 426574 65834 426658
rect 65254 426338 65426 426574
rect 65662 426338 65834 426574
rect 65254 390894 65834 426338
rect 65254 390658 65426 390894
rect 65662 390658 65834 390894
rect 65254 390574 65834 390658
rect 65254 390338 65426 390574
rect 65662 390338 65834 390574
rect 65254 354894 65834 390338
rect 65254 354658 65426 354894
rect 65662 354658 65834 354894
rect 65254 354574 65834 354658
rect 65254 354338 65426 354574
rect 65662 354338 65834 354574
rect 65254 318894 65834 354338
rect 65254 318658 65426 318894
rect 65662 318658 65834 318894
rect 65254 318574 65834 318658
rect 65254 318338 65426 318574
rect 65662 318338 65834 318574
rect 65254 282894 65834 318338
rect 65254 282658 65426 282894
rect 65662 282658 65834 282894
rect 65254 282574 65834 282658
rect 65254 282338 65426 282574
rect 65662 282338 65834 282574
rect 65254 246894 65834 282338
rect 65254 246658 65426 246894
rect 65662 246658 65834 246894
rect 65254 246574 65834 246658
rect 65254 246338 65426 246574
rect 65662 246338 65834 246574
rect 65254 210894 65834 246338
rect 65254 210658 65426 210894
rect 65662 210658 65834 210894
rect 65254 210574 65834 210658
rect 65254 210338 65426 210574
rect 65662 210338 65834 210574
rect 65254 174894 65834 210338
rect 65254 174658 65426 174894
rect 65662 174658 65834 174894
rect 65254 174574 65834 174658
rect 65254 174338 65426 174574
rect 65662 174338 65834 174574
rect 65254 138894 65834 174338
rect 65254 138658 65426 138894
rect 65662 138658 65834 138894
rect 65254 138574 65834 138658
rect 65254 138338 65426 138574
rect 65662 138338 65834 138574
rect 65254 102894 65834 138338
rect 65254 102658 65426 102894
rect 65662 102658 65834 102894
rect 65254 102574 65834 102658
rect 65254 102338 65426 102574
rect 65662 102338 65834 102574
rect 65254 66894 65834 102338
rect 65254 66658 65426 66894
rect 65662 66658 65834 66894
rect 65254 66574 65834 66658
rect 65254 66338 65426 66574
rect 65662 66338 65834 66574
rect 65254 30894 65834 66338
rect 65254 30658 65426 30894
rect 65662 30658 65834 30894
rect 65254 30574 65834 30658
rect 65254 30338 65426 30574
rect 65662 30338 65834 30574
rect 47254 -6102 47426 -5866
rect 47662 -6102 47834 -5866
rect 47254 -6186 47834 -6102
rect 47254 -6422 47426 -6186
rect 47662 -6422 47834 -6186
rect 47254 -7354 47834 -6422
rect 65254 -6786 65834 30338
rect 72814 704838 73394 705770
rect 72814 704602 72986 704838
rect 73222 704602 73394 704838
rect 72814 704518 73394 704602
rect 72814 704282 72986 704518
rect 73222 704282 73394 704518
rect 72814 686454 73394 704282
rect 72814 686218 72986 686454
rect 73222 686218 73394 686454
rect 72814 686134 73394 686218
rect 72814 685898 72986 686134
rect 73222 685898 73394 686134
rect 72814 650454 73394 685898
rect 72814 650218 72986 650454
rect 73222 650218 73394 650454
rect 72814 650134 73394 650218
rect 72814 649898 72986 650134
rect 73222 649898 73394 650134
rect 72814 614454 73394 649898
rect 72814 614218 72986 614454
rect 73222 614218 73394 614454
rect 72814 614134 73394 614218
rect 72814 613898 72986 614134
rect 73222 613898 73394 614134
rect 72814 578454 73394 613898
rect 72814 578218 72986 578454
rect 73222 578218 73394 578454
rect 72814 578134 73394 578218
rect 72814 577898 72986 578134
rect 73222 577898 73394 578134
rect 72814 542454 73394 577898
rect 72814 542218 72986 542454
rect 73222 542218 73394 542454
rect 72814 542134 73394 542218
rect 72814 541898 72986 542134
rect 73222 541898 73394 542134
rect 72814 506454 73394 541898
rect 72814 506218 72986 506454
rect 73222 506218 73394 506454
rect 72814 506134 73394 506218
rect 72814 505898 72986 506134
rect 73222 505898 73394 506134
rect 72814 470454 73394 505898
rect 72814 470218 72986 470454
rect 73222 470218 73394 470454
rect 72814 470134 73394 470218
rect 72814 469898 72986 470134
rect 73222 469898 73394 470134
rect 72814 434454 73394 469898
rect 72814 434218 72986 434454
rect 73222 434218 73394 434454
rect 72814 434134 73394 434218
rect 72814 433898 72986 434134
rect 73222 433898 73394 434134
rect 72814 398454 73394 433898
rect 72814 398218 72986 398454
rect 73222 398218 73394 398454
rect 72814 398134 73394 398218
rect 72814 397898 72986 398134
rect 73222 397898 73394 398134
rect 72814 362454 73394 397898
rect 72814 362218 72986 362454
rect 73222 362218 73394 362454
rect 72814 362134 73394 362218
rect 72814 361898 72986 362134
rect 73222 361898 73394 362134
rect 72814 326454 73394 361898
rect 72814 326218 72986 326454
rect 73222 326218 73394 326454
rect 72814 326134 73394 326218
rect 72814 325898 72986 326134
rect 73222 325898 73394 326134
rect 72814 290454 73394 325898
rect 72814 290218 72986 290454
rect 73222 290218 73394 290454
rect 72814 290134 73394 290218
rect 72814 289898 72986 290134
rect 73222 289898 73394 290134
rect 72814 254454 73394 289898
rect 72814 254218 72986 254454
rect 73222 254218 73394 254454
rect 72814 254134 73394 254218
rect 72814 253898 72986 254134
rect 73222 253898 73394 254134
rect 72814 218454 73394 253898
rect 72814 218218 72986 218454
rect 73222 218218 73394 218454
rect 72814 218134 73394 218218
rect 72814 217898 72986 218134
rect 73222 217898 73394 218134
rect 72814 182454 73394 217898
rect 72814 182218 72986 182454
rect 73222 182218 73394 182454
rect 72814 182134 73394 182218
rect 72814 181898 72986 182134
rect 73222 181898 73394 182134
rect 72814 146454 73394 181898
rect 72814 146218 72986 146454
rect 73222 146218 73394 146454
rect 72814 146134 73394 146218
rect 72814 145898 72986 146134
rect 73222 145898 73394 146134
rect 72814 110454 73394 145898
rect 72814 110218 72986 110454
rect 73222 110218 73394 110454
rect 72814 110134 73394 110218
rect 72814 109898 72986 110134
rect 73222 109898 73394 110134
rect 72814 74454 73394 109898
rect 72814 74218 72986 74454
rect 73222 74218 73394 74454
rect 72814 74134 73394 74218
rect 72814 73898 72986 74134
rect 73222 73898 73394 74134
rect 72814 38454 73394 73898
rect 72814 38218 72986 38454
rect 73222 38218 73394 38454
rect 72814 38134 73394 38218
rect 72814 37898 72986 38134
rect 73222 37898 73394 38134
rect 72814 2454 73394 37898
rect 72814 2218 72986 2454
rect 73222 2218 73394 2454
rect 72814 2134 73394 2218
rect 72814 1898 72986 2134
rect 73222 1898 73394 2134
rect 72814 -346 73394 1898
rect 72814 -582 72986 -346
rect 73222 -582 73394 -346
rect 72814 -666 73394 -582
rect 72814 -902 72986 -666
rect 73222 -902 73394 -666
rect 72814 -1834 73394 -902
rect 76294 689934 76874 706122
rect 76294 689698 76466 689934
rect 76702 689698 76874 689934
rect 76294 689614 76874 689698
rect 76294 689378 76466 689614
rect 76702 689378 76874 689614
rect 76294 653934 76874 689378
rect 76294 653698 76466 653934
rect 76702 653698 76874 653934
rect 76294 653614 76874 653698
rect 76294 653378 76466 653614
rect 76702 653378 76874 653614
rect 76294 617934 76874 653378
rect 76294 617698 76466 617934
rect 76702 617698 76874 617934
rect 76294 617614 76874 617698
rect 76294 617378 76466 617614
rect 76702 617378 76874 617614
rect 76294 581934 76874 617378
rect 76294 581698 76466 581934
rect 76702 581698 76874 581934
rect 76294 581614 76874 581698
rect 76294 581378 76466 581614
rect 76702 581378 76874 581614
rect 76294 545934 76874 581378
rect 76294 545698 76466 545934
rect 76702 545698 76874 545934
rect 76294 545614 76874 545698
rect 76294 545378 76466 545614
rect 76702 545378 76874 545614
rect 76294 509934 76874 545378
rect 76294 509698 76466 509934
rect 76702 509698 76874 509934
rect 76294 509614 76874 509698
rect 76294 509378 76466 509614
rect 76702 509378 76874 509614
rect 76294 473934 76874 509378
rect 76294 473698 76466 473934
rect 76702 473698 76874 473934
rect 76294 473614 76874 473698
rect 76294 473378 76466 473614
rect 76702 473378 76874 473614
rect 76294 437934 76874 473378
rect 76294 437698 76466 437934
rect 76702 437698 76874 437934
rect 76294 437614 76874 437698
rect 76294 437378 76466 437614
rect 76702 437378 76874 437614
rect 76294 401934 76874 437378
rect 76294 401698 76466 401934
rect 76702 401698 76874 401934
rect 76294 401614 76874 401698
rect 76294 401378 76466 401614
rect 76702 401378 76874 401614
rect 76294 365934 76874 401378
rect 76294 365698 76466 365934
rect 76702 365698 76874 365934
rect 76294 365614 76874 365698
rect 76294 365378 76466 365614
rect 76702 365378 76874 365614
rect 76294 329934 76874 365378
rect 76294 329698 76466 329934
rect 76702 329698 76874 329934
rect 76294 329614 76874 329698
rect 76294 329378 76466 329614
rect 76702 329378 76874 329614
rect 76294 293934 76874 329378
rect 76294 293698 76466 293934
rect 76702 293698 76874 293934
rect 76294 293614 76874 293698
rect 76294 293378 76466 293614
rect 76702 293378 76874 293614
rect 76294 257934 76874 293378
rect 76294 257698 76466 257934
rect 76702 257698 76874 257934
rect 76294 257614 76874 257698
rect 76294 257378 76466 257614
rect 76702 257378 76874 257614
rect 76294 221934 76874 257378
rect 76294 221698 76466 221934
rect 76702 221698 76874 221934
rect 76294 221614 76874 221698
rect 76294 221378 76466 221614
rect 76702 221378 76874 221614
rect 76294 185934 76874 221378
rect 76294 185698 76466 185934
rect 76702 185698 76874 185934
rect 76294 185614 76874 185698
rect 76294 185378 76466 185614
rect 76702 185378 76874 185614
rect 76294 149934 76874 185378
rect 76294 149698 76466 149934
rect 76702 149698 76874 149934
rect 76294 149614 76874 149698
rect 76294 149378 76466 149614
rect 76702 149378 76874 149614
rect 76294 113934 76874 149378
rect 76294 113698 76466 113934
rect 76702 113698 76874 113934
rect 76294 113614 76874 113698
rect 76294 113378 76466 113614
rect 76702 113378 76874 113614
rect 76294 77934 76874 113378
rect 76294 77698 76466 77934
rect 76702 77698 76874 77934
rect 76294 77614 76874 77698
rect 76294 77378 76466 77614
rect 76702 77378 76874 77614
rect 76294 41934 76874 77378
rect 76294 41698 76466 41934
rect 76702 41698 76874 41934
rect 76294 41614 76874 41698
rect 76294 41378 76466 41614
rect 76702 41378 76874 41614
rect 76294 5934 76874 41378
rect 76294 5698 76466 5934
rect 76702 5698 76874 5934
rect 76294 5614 76874 5698
rect 76294 5378 76466 5614
rect 76702 5378 76874 5614
rect 76294 -2186 76874 5378
rect 76294 -2422 76466 -2186
rect 76702 -2422 76874 -2186
rect 76294 -2506 76874 -2422
rect 76294 -2742 76466 -2506
rect 76702 -2742 76874 -2506
rect 76294 -3674 76874 -2742
rect 79774 693414 80354 707962
rect 79774 693178 79946 693414
rect 80182 693178 80354 693414
rect 79774 693094 80354 693178
rect 79774 692858 79946 693094
rect 80182 692858 80354 693094
rect 79774 657414 80354 692858
rect 79774 657178 79946 657414
rect 80182 657178 80354 657414
rect 79774 657094 80354 657178
rect 79774 656858 79946 657094
rect 80182 656858 80354 657094
rect 79774 621414 80354 656858
rect 79774 621178 79946 621414
rect 80182 621178 80354 621414
rect 79774 621094 80354 621178
rect 79774 620858 79946 621094
rect 80182 620858 80354 621094
rect 79774 585414 80354 620858
rect 79774 585178 79946 585414
rect 80182 585178 80354 585414
rect 79774 585094 80354 585178
rect 79774 584858 79946 585094
rect 80182 584858 80354 585094
rect 79774 549414 80354 584858
rect 79774 549178 79946 549414
rect 80182 549178 80354 549414
rect 79774 549094 80354 549178
rect 79774 548858 79946 549094
rect 80182 548858 80354 549094
rect 79774 513414 80354 548858
rect 79774 513178 79946 513414
rect 80182 513178 80354 513414
rect 79774 513094 80354 513178
rect 79774 512858 79946 513094
rect 80182 512858 80354 513094
rect 79774 477414 80354 512858
rect 79774 477178 79946 477414
rect 80182 477178 80354 477414
rect 79774 477094 80354 477178
rect 79774 476858 79946 477094
rect 80182 476858 80354 477094
rect 79774 441414 80354 476858
rect 79774 441178 79946 441414
rect 80182 441178 80354 441414
rect 79774 441094 80354 441178
rect 79774 440858 79946 441094
rect 80182 440858 80354 441094
rect 79774 405414 80354 440858
rect 79774 405178 79946 405414
rect 80182 405178 80354 405414
rect 79774 405094 80354 405178
rect 79774 404858 79946 405094
rect 80182 404858 80354 405094
rect 79774 369414 80354 404858
rect 79774 369178 79946 369414
rect 80182 369178 80354 369414
rect 79774 369094 80354 369178
rect 79774 368858 79946 369094
rect 80182 368858 80354 369094
rect 79774 333414 80354 368858
rect 79774 333178 79946 333414
rect 80182 333178 80354 333414
rect 79774 333094 80354 333178
rect 79774 332858 79946 333094
rect 80182 332858 80354 333094
rect 79774 297414 80354 332858
rect 79774 297178 79946 297414
rect 80182 297178 80354 297414
rect 79774 297094 80354 297178
rect 79774 296858 79946 297094
rect 80182 296858 80354 297094
rect 79774 261414 80354 296858
rect 79774 261178 79946 261414
rect 80182 261178 80354 261414
rect 79774 261094 80354 261178
rect 79774 260858 79946 261094
rect 80182 260858 80354 261094
rect 79774 225414 80354 260858
rect 79774 225178 79946 225414
rect 80182 225178 80354 225414
rect 79774 225094 80354 225178
rect 79774 224858 79946 225094
rect 80182 224858 80354 225094
rect 79774 189414 80354 224858
rect 79774 189178 79946 189414
rect 80182 189178 80354 189414
rect 79774 189094 80354 189178
rect 79774 188858 79946 189094
rect 80182 188858 80354 189094
rect 79774 153414 80354 188858
rect 79774 153178 79946 153414
rect 80182 153178 80354 153414
rect 79774 153094 80354 153178
rect 79774 152858 79946 153094
rect 80182 152858 80354 153094
rect 79774 117414 80354 152858
rect 79774 117178 79946 117414
rect 80182 117178 80354 117414
rect 79774 117094 80354 117178
rect 79774 116858 79946 117094
rect 80182 116858 80354 117094
rect 79774 81414 80354 116858
rect 79774 81178 79946 81414
rect 80182 81178 80354 81414
rect 79774 81094 80354 81178
rect 79774 80858 79946 81094
rect 80182 80858 80354 81094
rect 79774 45414 80354 80858
rect 79774 45178 79946 45414
rect 80182 45178 80354 45414
rect 79774 45094 80354 45178
rect 79774 44858 79946 45094
rect 80182 44858 80354 45094
rect 79774 9414 80354 44858
rect 79774 9178 79946 9414
rect 80182 9178 80354 9414
rect 79774 9094 80354 9178
rect 79774 8858 79946 9094
rect 80182 8858 80354 9094
rect 79774 -4026 80354 8858
rect 79774 -4262 79946 -4026
rect 80182 -4262 80354 -4026
rect 79774 -4346 80354 -4262
rect 79774 -4582 79946 -4346
rect 80182 -4582 80354 -4346
rect 79774 -5514 80354 -4582
rect 83254 696894 83834 709802
rect 101254 711278 101834 711290
rect 101254 711042 101426 711278
rect 101662 711042 101834 711278
rect 101254 710958 101834 711042
rect 101254 710722 101426 710958
rect 101662 710722 101834 710958
rect 97774 709438 98354 709450
rect 97774 709202 97946 709438
rect 98182 709202 98354 709438
rect 97774 709118 98354 709202
rect 97774 708882 97946 709118
rect 98182 708882 98354 709118
rect 94294 707598 94874 707610
rect 94294 707362 94466 707598
rect 94702 707362 94874 707598
rect 94294 707278 94874 707362
rect 94294 707042 94466 707278
rect 94702 707042 94874 707278
rect 83254 696658 83426 696894
rect 83662 696658 83834 696894
rect 83254 696574 83834 696658
rect 83254 696338 83426 696574
rect 83662 696338 83834 696574
rect 83254 660894 83834 696338
rect 83254 660658 83426 660894
rect 83662 660658 83834 660894
rect 83254 660574 83834 660658
rect 83254 660338 83426 660574
rect 83662 660338 83834 660574
rect 83254 624894 83834 660338
rect 83254 624658 83426 624894
rect 83662 624658 83834 624894
rect 83254 624574 83834 624658
rect 83254 624338 83426 624574
rect 83662 624338 83834 624574
rect 83254 588894 83834 624338
rect 83254 588658 83426 588894
rect 83662 588658 83834 588894
rect 83254 588574 83834 588658
rect 83254 588338 83426 588574
rect 83662 588338 83834 588574
rect 83254 552894 83834 588338
rect 83254 552658 83426 552894
rect 83662 552658 83834 552894
rect 83254 552574 83834 552658
rect 83254 552338 83426 552574
rect 83662 552338 83834 552574
rect 83254 516894 83834 552338
rect 83254 516658 83426 516894
rect 83662 516658 83834 516894
rect 83254 516574 83834 516658
rect 83254 516338 83426 516574
rect 83662 516338 83834 516574
rect 83254 480894 83834 516338
rect 83254 480658 83426 480894
rect 83662 480658 83834 480894
rect 83254 480574 83834 480658
rect 83254 480338 83426 480574
rect 83662 480338 83834 480574
rect 83254 444894 83834 480338
rect 83254 444658 83426 444894
rect 83662 444658 83834 444894
rect 83254 444574 83834 444658
rect 83254 444338 83426 444574
rect 83662 444338 83834 444574
rect 83254 408894 83834 444338
rect 83254 408658 83426 408894
rect 83662 408658 83834 408894
rect 83254 408574 83834 408658
rect 83254 408338 83426 408574
rect 83662 408338 83834 408574
rect 83254 372894 83834 408338
rect 83254 372658 83426 372894
rect 83662 372658 83834 372894
rect 83254 372574 83834 372658
rect 83254 372338 83426 372574
rect 83662 372338 83834 372574
rect 83254 336894 83834 372338
rect 83254 336658 83426 336894
rect 83662 336658 83834 336894
rect 83254 336574 83834 336658
rect 83254 336338 83426 336574
rect 83662 336338 83834 336574
rect 83254 300894 83834 336338
rect 83254 300658 83426 300894
rect 83662 300658 83834 300894
rect 83254 300574 83834 300658
rect 83254 300338 83426 300574
rect 83662 300338 83834 300574
rect 83254 264894 83834 300338
rect 83254 264658 83426 264894
rect 83662 264658 83834 264894
rect 83254 264574 83834 264658
rect 83254 264338 83426 264574
rect 83662 264338 83834 264574
rect 83254 228894 83834 264338
rect 83254 228658 83426 228894
rect 83662 228658 83834 228894
rect 83254 228574 83834 228658
rect 83254 228338 83426 228574
rect 83662 228338 83834 228574
rect 83254 192894 83834 228338
rect 83254 192658 83426 192894
rect 83662 192658 83834 192894
rect 83254 192574 83834 192658
rect 83254 192338 83426 192574
rect 83662 192338 83834 192574
rect 83254 156894 83834 192338
rect 83254 156658 83426 156894
rect 83662 156658 83834 156894
rect 83254 156574 83834 156658
rect 83254 156338 83426 156574
rect 83662 156338 83834 156574
rect 83254 120894 83834 156338
rect 83254 120658 83426 120894
rect 83662 120658 83834 120894
rect 83254 120574 83834 120658
rect 83254 120338 83426 120574
rect 83662 120338 83834 120574
rect 83254 84894 83834 120338
rect 83254 84658 83426 84894
rect 83662 84658 83834 84894
rect 83254 84574 83834 84658
rect 83254 84338 83426 84574
rect 83662 84338 83834 84574
rect 83254 48894 83834 84338
rect 83254 48658 83426 48894
rect 83662 48658 83834 48894
rect 83254 48574 83834 48658
rect 83254 48338 83426 48574
rect 83662 48338 83834 48574
rect 83254 12894 83834 48338
rect 83254 12658 83426 12894
rect 83662 12658 83834 12894
rect 83254 12574 83834 12658
rect 83254 12338 83426 12574
rect 83662 12338 83834 12574
rect 65254 -7022 65426 -6786
rect 65662 -7022 65834 -6786
rect 65254 -7106 65834 -7022
rect 65254 -7342 65426 -7106
rect 65662 -7342 65834 -7106
rect 65254 -7354 65834 -7342
rect 83254 -5866 83834 12338
rect 90814 705758 91394 705770
rect 90814 705522 90986 705758
rect 91222 705522 91394 705758
rect 90814 705438 91394 705522
rect 90814 705202 90986 705438
rect 91222 705202 91394 705438
rect 90814 668454 91394 705202
rect 90814 668218 90986 668454
rect 91222 668218 91394 668454
rect 90814 668134 91394 668218
rect 90814 667898 90986 668134
rect 91222 667898 91394 668134
rect 90814 632454 91394 667898
rect 90814 632218 90986 632454
rect 91222 632218 91394 632454
rect 90814 632134 91394 632218
rect 90814 631898 90986 632134
rect 91222 631898 91394 632134
rect 90814 596454 91394 631898
rect 90814 596218 90986 596454
rect 91222 596218 91394 596454
rect 90814 596134 91394 596218
rect 90814 595898 90986 596134
rect 91222 595898 91394 596134
rect 90814 560454 91394 595898
rect 90814 560218 90986 560454
rect 91222 560218 91394 560454
rect 90814 560134 91394 560218
rect 90814 559898 90986 560134
rect 91222 559898 91394 560134
rect 90814 524454 91394 559898
rect 90814 524218 90986 524454
rect 91222 524218 91394 524454
rect 90814 524134 91394 524218
rect 90814 523898 90986 524134
rect 91222 523898 91394 524134
rect 90814 488454 91394 523898
rect 90814 488218 90986 488454
rect 91222 488218 91394 488454
rect 90814 488134 91394 488218
rect 90814 487898 90986 488134
rect 91222 487898 91394 488134
rect 90814 452454 91394 487898
rect 90814 452218 90986 452454
rect 91222 452218 91394 452454
rect 90814 452134 91394 452218
rect 90814 451898 90986 452134
rect 91222 451898 91394 452134
rect 90814 416454 91394 451898
rect 90814 416218 90986 416454
rect 91222 416218 91394 416454
rect 90814 416134 91394 416218
rect 90814 415898 90986 416134
rect 91222 415898 91394 416134
rect 90814 380454 91394 415898
rect 90814 380218 90986 380454
rect 91222 380218 91394 380454
rect 90814 380134 91394 380218
rect 90814 379898 90986 380134
rect 91222 379898 91394 380134
rect 90814 344454 91394 379898
rect 90814 344218 90986 344454
rect 91222 344218 91394 344454
rect 90814 344134 91394 344218
rect 90814 343898 90986 344134
rect 91222 343898 91394 344134
rect 90814 308454 91394 343898
rect 90814 308218 90986 308454
rect 91222 308218 91394 308454
rect 90814 308134 91394 308218
rect 90814 307898 90986 308134
rect 91222 307898 91394 308134
rect 90814 272454 91394 307898
rect 90814 272218 90986 272454
rect 91222 272218 91394 272454
rect 90814 272134 91394 272218
rect 90814 271898 90986 272134
rect 91222 271898 91394 272134
rect 90814 236454 91394 271898
rect 90814 236218 90986 236454
rect 91222 236218 91394 236454
rect 90814 236134 91394 236218
rect 90814 235898 90986 236134
rect 91222 235898 91394 236134
rect 90814 200454 91394 235898
rect 90814 200218 90986 200454
rect 91222 200218 91394 200454
rect 90814 200134 91394 200218
rect 90814 199898 90986 200134
rect 91222 199898 91394 200134
rect 90814 164454 91394 199898
rect 90814 164218 90986 164454
rect 91222 164218 91394 164454
rect 90814 164134 91394 164218
rect 90814 163898 90986 164134
rect 91222 163898 91394 164134
rect 90814 128454 91394 163898
rect 90814 128218 90986 128454
rect 91222 128218 91394 128454
rect 90814 128134 91394 128218
rect 90814 127898 90986 128134
rect 91222 127898 91394 128134
rect 90814 92454 91394 127898
rect 90814 92218 90986 92454
rect 91222 92218 91394 92454
rect 90814 92134 91394 92218
rect 90814 91898 90986 92134
rect 91222 91898 91394 92134
rect 90814 56454 91394 91898
rect 90814 56218 90986 56454
rect 91222 56218 91394 56454
rect 90814 56134 91394 56218
rect 90814 55898 90986 56134
rect 91222 55898 91394 56134
rect 90814 20454 91394 55898
rect 90814 20218 90986 20454
rect 91222 20218 91394 20454
rect 90814 20134 91394 20218
rect 90814 19898 90986 20134
rect 91222 19898 91394 20134
rect 90814 -1266 91394 19898
rect 90814 -1502 90986 -1266
rect 91222 -1502 91394 -1266
rect 90814 -1586 91394 -1502
rect 90814 -1822 90986 -1586
rect 91222 -1822 91394 -1586
rect 90814 -1834 91394 -1822
rect 94294 671934 94874 707042
rect 94294 671698 94466 671934
rect 94702 671698 94874 671934
rect 94294 671614 94874 671698
rect 94294 671378 94466 671614
rect 94702 671378 94874 671614
rect 94294 635934 94874 671378
rect 94294 635698 94466 635934
rect 94702 635698 94874 635934
rect 94294 635614 94874 635698
rect 94294 635378 94466 635614
rect 94702 635378 94874 635614
rect 94294 599934 94874 635378
rect 94294 599698 94466 599934
rect 94702 599698 94874 599934
rect 94294 599614 94874 599698
rect 94294 599378 94466 599614
rect 94702 599378 94874 599614
rect 94294 563934 94874 599378
rect 94294 563698 94466 563934
rect 94702 563698 94874 563934
rect 94294 563614 94874 563698
rect 94294 563378 94466 563614
rect 94702 563378 94874 563614
rect 94294 527934 94874 563378
rect 94294 527698 94466 527934
rect 94702 527698 94874 527934
rect 94294 527614 94874 527698
rect 94294 527378 94466 527614
rect 94702 527378 94874 527614
rect 94294 491934 94874 527378
rect 94294 491698 94466 491934
rect 94702 491698 94874 491934
rect 94294 491614 94874 491698
rect 94294 491378 94466 491614
rect 94702 491378 94874 491614
rect 94294 455934 94874 491378
rect 94294 455698 94466 455934
rect 94702 455698 94874 455934
rect 94294 455614 94874 455698
rect 94294 455378 94466 455614
rect 94702 455378 94874 455614
rect 94294 419934 94874 455378
rect 94294 419698 94466 419934
rect 94702 419698 94874 419934
rect 94294 419614 94874 419698
rect 94294 419378 94466 419614
rect 94702 419378 94874 419614
rect 94294 383934 94874 419378
rect 94294 383698 94466 383934
rect 94702 383698 94874 383934
rect 94294 383614 94874 383698
rect 94294 383378 94466 383614
rect 94702 383378 94874 383614
rect 94294 347934 94874 383378
rect 94294 347698 94466 347934
rect 94702 347698 94874 347934
rect 94294 347614 94874 347698
rect 94294 347378 94466 347614
rect 94702 347378 94874 347614
rect 94294 311934 94874 347378
rect 94294 311698 94466 311934
rect 94702 311698 94874 311934
rect 94294 311614 94874 311698
rect 94294 311378 94466 311614
rect 94702 311378 94874 311614
rect 94294 275934 94874 311378
rect 94294 275698 94466 275934
rect 94702 275698 94874 275934
rect 94294 275614 94874 275698
rect 94294 275378 94466 275614
rect 94702 275378 94874 275614
rect 94294 239934 94874 275378
rect 94294 239698 94466 239934
rect 94702 239698 94874 239934
rect 94294 239614 94874 239698
rect 94294 239378 94466 239614
rect 94702 239378 94874 239614
rect 94294 203934 94874 239378
rect 94294 203698 94466 203934
rect 94702 203698 94874 203934
rect 94294 203614 94874 203698
rect 94294 203378 94466 203614
rect 94702 203378 94874 203614
rect 94294 167934 94874 203378
rect 94294 167698 94466 167934
rect 94702 167698 94874 167934
rect 94294 167614 94874 167698
rect 94294 167378 94466 167614
rect 94702 167378 94874 167614
rect 94294 131934 94874 167378
rect 94294 131698 94466 131934
rect 94702 131698 94874 131934
rect 94294 131614 94874 131698
rect 94294 131378 94466 131614
rect 94702 131378 94874 131614
rect 94294 95934 94874 131378
rect 94294 95698 94466 95934
rect 94702 95698 94874 95934
rect 94294 95614 94874 95698
rect 94294 95378 94466 95614
rect 94702 95378 94874 95614
rect 94294 59934 94874 95378
rect 94294 59698 94466 59934
rect 94702 59698 94874 59934
rect 94294 59614 94874 59698
rect 94294 59378 94466 59614
rect 94702 59378 94874 59614
rect 94294 23934 94874 59378
rect 94294 23698 94466 23934
rect 94702 23698 94874 23934
rect 94294 23614 94874 23698
rect 94294 23378 94466 23614
rect 94702 23378 94874 23614
rect 94294 -3106 94874 23378
rect 94294 -3342 94466 -3106
rect 94702 -3342 94874 -3106
rect 94294 -3426 94874 -3342
rect 94294 -3662 94466 -3426
rect 94702 -3662 94874 -3426
rect 94294 -3674 94874 -3662
rect 97774 675414 98354 708882
rect 97774 675178 97946 675414
rect 98182 675178 98354 675414
rect 97774 675094 98354 675178
rect 97774 674858 97946 675094
rect 98182 674858 98354 675094
rect 97774 639414 98354 674858
rect 97774 639178 97946 639414
rect 98182 639178 98354 639414
rect 97774 639094 98354 639178
rect 97774 638858 97946 639094
rect 98182 638858 98354 639094
rect 97774 603414 98354 638858
rect 97774 603178 97946 603414
rect 98182 603178 98354 603414
rect 97774 603094 98354 603178
rect 97774 602858 97946 603094
rect 98182 602858 98354 603094
rect 97774 567414 98354 602858
rect 97774 567178 97946 567414
rect 98182 567178 98354 567414
rect 97774 567094 98354 567178
rect 97774 566858 97946 567094
rect 98182 566858 98354 567094
rect 97774 531414 98354 566858
rect 97774 531178 97946 531414
rect 98182 531178 98354 531414
rect 97774 531094 98354 531178
rect 97774 530858 97946 531094
rect 98182 530858 98354 531094
rect 97774 495414 98354 530858
rect 97774 495178 97946 495414
rect 98182 495178 98354 495414
rect 97774 495094 98354 495178
rect 97774 494858 97946 495094
rect 98182 494858 98354 495094
rect 97774 459414 98354 494858
rect 97774 459178 97946 459414
rect 98182 459178 98354 459414
rect 97774 459094 98354 459178
rect 97774 458858 97946 459094
rect 98182 458858 98354 459094
rect 97774 423414 98354 458858
rect 97774 423178 97946 423414
rect 98182 423178 98354 423414
rect 97774 423094 98354 423178
rect 97774 422858 97946 423094
rect 98182 422858 98354 423094
rect 97774 387414 98354 422858
rect 97774 387178 97946 387414
rect 98182 387178 98354 387414
rect 97774 387094 98354 387178
rect 97774 386858 97946 387094
rect 98182 386858 98354 387094
rect 97774 351414 98354 386858
rect 97774 351178 97946 351414
rect 98182 351178 98354 351414
rect 97774 351094 98354 351178
rect 97774 350858 97946 351094
rect 98182 350858 98354 351094
rect 97774 315414 98354 350858
rect 97774 315178 97946 315414
rect 98182 315178 98354 315414
rect 97774 315094 98354 315178
rect 97774 314858 97946 315094
rect 98182 314858 98354 315094
rect 97774 279414 98354 314858
rect 97774 279178 97946 279414
rect 98182 279178 98354 279414
rect 97774 279094 98354 279178
rect 97774 278858 97946 279094
rect 98182 278858 98354 279094
rect 97774 243414 98354 278858
rect 97774 243178 97946 243414
rect 98182 243178 98354 243414
rect 97774 243094 98354 243178
rect 97774 242858 97946 243094
rect 98182 242858 98354 243094
rect 97774 207414 98354 242858
rect 97774 207178 97946 207414
rect 98182 207178 98354 207414
rect 97774 207094 98354 207178
rect 97774 206858 97946 207094
rect 98182 206858 98354 207094
rect 97774 171414 98354 206858
rect 97774 171178 97946 171414
rect 98182 171178 98354 171414
rect 97774 171094 98354 171178
rect 97774 170858 97946 171094
rect 98182 170858 98354 171094
rect 97774 135414 98354 170858
rect 97774 135178 97946 135414
rect 98182 135178 98354 135414
rect 97774 135094 98354 135178
rect 97774 134858 97946 135094
rect 98182 134858 98354 135094
rect 97774 99414 98354 134858
rect 97774 99178 97946 99414
rect 98182 99178 98354 99414
rect 97774 99094 98354 99178
rect 97774 98858 97946 99094
rect 98182 98858 98354 99094
rect 97774 63414 98354 98858
rect 97774 63178 97946 63414
rect 98182 63178 98354 63414
rect 97774 63094 98354 63178
rect 97774 62858 97946 63094
rect 98182 62858 98354 63094
rect 97774 27414 98354 62858
rect 97774 27178 97946 27414
rect 98182 27178 98354 27414
rect 97774 27094 98354 27178
rect 97774 26858 97946 27094
rect 98182 26858 98354 27094
rect 97774 -4946 98354 26858
rect 97774 -5182 97946 -4946
rect 98182 -5182 98354 -4946
rect 97774 -5266 98354 -5182
rect 97774 -5502 97946 -5266
rect 98182 -5502 98354 -5266
rect 97774 -5514 98354 -5502
rect 101254 678894 101834 710722
rect 119254 710358 119834 711290
rect 119254 710122 119426 710358
rect 119662 710122 119834 710358
rect 119254 710038 119834 710122
rect 119254 709802 119426 710038
rect 119662 709802 119834 710038
rect 115774 708518 116354 709450
rect 115774 708282 115946 708518
rect 116182 708282 116354 708518
rect 115774 708198 116354 708282
rect 115774 707962 115946 708198
rect 116182 707962 116354 708198
rect 112294 706678 112874 707610
rect 112294 706442 112466 706678
rect 112702 706442 112874 706678
rect 112294 706358 112874 706442
rect 112294 706122 112466 706358
rect 112702 706122 112874 706358
rect 101254 678658 101426 678894
rect 101662 678658 101834 678894
rect 101254 678574 101834 678658
rect 101254 678338 101426 678574
rect 101662 678338 101834 678574
rect 101254 642894 101834 678338
rect 101254 642658 101426 642894
rect 101662 642658 101834 642894
rect 101254 642574 101834 642658
rect 101254 642338 101426 642574
rect 101662 642338 101834 642574
rect 101254 606894 101834 642338
rect 101254 606658 101426 606894
rect 101662 606658 101834 606894
rect 101254 606574 101834 606658
rect 101254 606338 101426 606574
rect 101662 606338 101834 606574
rect 101254 570894 101834 606338
rect 101254 570658 101426 570894
rect 101662 570658 101834 570894
rect 101254 570574 101834 570658
rect 101254 570338 101426 570574
rect 101662 570338 101834 570574
rect 101254 534894 101834 570338
rect 101254 534658 101426 534894
rect 101662 534658 101834 534894
rect 101254 534574 101834 534658
rect 101254 534338 101426 534574
rect 101662 534338 101834 534574
rect 101254 498894 101834 534338
rect 101254 498658 101426 498894
rect 101662 498658 101834 498894
rect 101254 498574 101834 498658
rect 101254 498338 101426 498574
rect 101662 498338 101834 498574
rect 101254 462894 101834 498338
rect 101254 462658 101426 462894
rect 101662 462658 101834 462894
rect 101254 462574 101834 462658
rect 101254 462338 101426 462574
rect 101662 462338 101834 462574
rect 101254 426894 101834 462338
rect 101254 426658 101426 426894
rect 101662 426658 101834 426894
rect 101254 426574 101834 426658
rect 101254 426338 101426 426574
rect 101662 426338 101834 426574
rect 101254 390894 101834 426338
rect 101254 390658 101426 390894
rect 101662 390658 101834 390894
rect 101254 390574 101834 390658
rect 101254 390338 101426 390574
rect 101662 390338 101834 390574
rect 101254 354894 101834 390338
rect 101254 354658 101426 354894
rect 101662 354658 101834 354894
rect 101254 354574 101834 354658
rect 101254 354338 101426 354574
rect 101662 354338 101834 354574
rect 101254 318894 101834 354338
rect 101254 318658 101426 318894
rect 101662 318658 101834 318894
rect 101254 318574 101834 318658
rect 101254 318338 101426 318574
rect 101662 318338 101834 318574
rect 101254 282894 101834 318338
rect 101254 282658 101426 282894
rect 101662 282658 101834 282894
rect 101254 282574 101834 282658
rect 101254 282338 101426 282574
rect 101662 282338 101834 282574
rect 101254 246894 101834 282338
rect 101254 246658 101426 246894
rect 101662 246658 101834 246894
rect 101254 246574 101834 246658
rect 101254 246338 101426 246574
rect 101662 246338 101834 246574
rect 101254 210894 101834 246338
rect 101254 210658 101426 210894
rect 101662 210658 101834 210894
rect 101254 210574 101834 210658
rect 101254 210338 101426 210574
rect 101662 210338 101834 210574
rect 101254 174894 101834 210338
rect 101254 174658 101426 174894
rect 101662 174658 101834 174894
rect 101254 174574 101834 174658
rect 101254 174338 101426 174574
rect 101662 174338 101834 174574
rect 101254 138894 101834 174338
rect 101254 138658 101426 138894
rect 101662 138658 101834 138894
rect 101254 138574 101834 138658
rect 101254 138338 101426 138574
rect 101662 138338 101834 138574
rect 101254 102894 101834 138338
rect 101254 102658 101426 102894
rect 101662 102658 101834 102894
rect 101254 102574 101834 102658
rect 101254 102338 101426 102574
rect 101662 102338 101834 102574
rect 101254 66894 101834 102338
rect 101254 66658 101426 66894
rect 101662 66658 101834 66894
rect 101254 66574 101834 66658
rect 101254 66338 101426 66574
rect 101662 66338 101834 66574
rect 101254 30894 101834 66338
rect 101254 30658 101426 30894
rect 101662 30658 101834 30894
rect 101254 30574 101834 30658
rect 101254 30338 101426 30574
rect 101662 30338 101834 30574
rect 83254 -6102 83426 -5866
rect 83662 -6102 83834 -5866
rect 83254 -6186 83834 -6102
rect 83254 -6422 83426 -6186
rect 83662 -6422 83834 -6186
rect 83254 -7354 83834 -6422
rect 101254 -6786 101834 30338
rect 108814 704838 109394 705770
rect 108814 704602 108986 704838
rect 109222 704602 109394 704838
rect 108814 704518 109394 704602
rect 108814 704282 108986 704518
rect 109222 704282 109394 704518
rect 108814 686454 109394 704282
rect 108814 686218 108986 686454
rect 109222 686218 109394 686454
rect 108814 686134 109394 686218
rect 108814 685898 108986 686134
rect 109222 685898 109394 686134
rect 108814 650454 109394 685898
rect 108814 650218 108986 650454
rect 109222 650218 109394 650454
rect 108814 650134 109394 650218
rect 108814 649898 108986 650134
rect 109222 649898 109394 650134
rect 108814 614454 109394 649898
rect 108814 614218 108986 614454
rect 109222 614218 109394 614454
rect 108814 614134 109394 614218
rect 108814 613898 108986 614134
rect 109222 613898 109394 614134
rect 108814 578454 109394 613898
rect 108814 578218 108986 578454
rect 109222 578218 109394 578454
rect 108814 578134 109394 578218
rect 108814 577898 108986 578134
rect 109222 577898 109394 578134
rect 108814 542454 109394 577898
rect 108814 542218 108986 542454
rect 109222 542218 109394 542454
rect 108814 542134 109394 542218
rect 108814 541898 108986 542134
rect 109222 541898 109394 542134
rect 108814 506454 109394 541898
rect 108814 506218 108986 506454
rect 109222 506218 109394 506454
rect 108814 506134 109394 506218
rect 108814 505898 108986 506134
rect 109222 505898 109394 506134
rect 108814 470454 109394 505898
rect 108814 470218 108986 470454
rect 109222 470218 109394 470454
rect 108814 470134 109394 470218
rect 108814 469898 108986 470134
rect 109222 469898 109394 470134
rect 108814 434454 109394 469898
rect 108814 434218 108986 434454
rect 109222 434218 109394 434454
rect 108814 434134 109394 434218
rect 108814 433898 108986 434134
rect 109222 433898 109394 434134
rect 108814 398454 109394 433898
rect 108814 398218 108986 398454
rect 109222 398218 109394 398454
rect 108814 398134 109394 398218
rect 108814 397898 108986 398134
rect 109222 397898 109394 398134
rect 108814 362454 109394 397898
rect 108814 362218 108986 362454
rect 109222 362218 109394 362454
rect 108814 362134 109394 362218
rect 108814 361898 108986 362134
rect 109222 361898 109394 362134
rect 108814 326454 109394 361898
rect 108814 326218 108986 326454
rect 109222 326218 109394 326454
rect 108814 326134 109394 326218
rect 108814 325898 108986 326134
rect 109222 325898 109394 326134
rect 108814 290454 109394 325898
rect 108814 290218 108986 290454
rect 109222 290218 109394 290454
rect 108814 290134 109394 290218
rect 108814 289898 108986 290134
rect 109222 289898 109394 290134
rect 108814 254454 109394 289898
rect 108814 254218 108986 254454
rect 109222 254218 109394 254454
rect 108814 254134 109394 254218
rect 108814 253898 108986 254134
rect 109222 253898 109394 254134
rect 108814 218454 109394 253898
rect 108814 218218 108986 218454
rect 109222 218218 109394 218454
rect 108814 218134 109394 218218
rect 108814 217898 108986 218134
rect 109222 217898 109394 218134
rect 108814 182454 109394 217898
rect 108814 182218 108986 182454
rect 109222 182218 109394 182454
rect 108814 182134 109394 182218
rect 108814 181898 108986 182134
rect 109222 181898 109394 182134
rect 108814 146454 109394 181898
rect 108814 146218 108986 146454
rect 109222 146218 109394 146454
rect 108814 146134 109394 146218
rect 108814 145898 108986 146134
rect 109222 145898 109394 146134
rect 108814 110454 109394 145898
rect 108814 110218 108986 110454
rect 109222 110218 109394 110454
rect 108814 110134 109394 110218
rect 108814 109898 108986 110134
rect 109222 109898 109394 110134
rect 108814 74454 109394 109898
rect 108814 74218 108986 74454
rect 109222 74218 109394 74454
rect 108814 74134 109394 74218
rect 108814 73898 108986 74134
rect 109222 73898 109394 74134
rect 108814 38454 109394 73898
rect 108814 38218 108986 38454
rect 109222 38218 109394 38454
rect 108814 38134 109394 38218
rect 108814 37898 108986 38134
rect 109222 37898 109394 38134
rect 108814 2454 109394 37898
rect 108814 2218 108986 2454
rect 109222 2218 109394 2454
rect 108814 2134 109394 2218
rect 108814 1898 108986 2134
rect 109222 1898 109394 2134
rect 108814 -346 109394 1898
rect 108814 -582 108986 -346
rect 109222 -582 109394 -346
rect 108814 -666 109394 -582
rect 108814 -902 108986 -666
rect 109222 -902 109394 -666
rect 108814 -1834 109394 -902
rect 112294 689934 112874 706122
rect 112294 689698 112466 689934
rect 112702 689698 112874 689934
rect 112294 689614 112874 689698
rect 112294 689378 112466 689614
rect 112702 689378 112874 689614
rect 112294 653934 112874 689378
rect 112294 653698 112466 653934
rect 112702 653698 112874 653934
rect 112294 653614 112874 653698
rect 112294 653378 112466 653614
rect 112702 653378 112874 653614
rect 112294 617934 112874 653378
rect 112294 617698 112466 617934
rect 112702 617698 112874 617934
rect 112294 617614 112874 617698
rect 112294 617378 112466 617614
rect 112702 617378 112874 617614
rect 112294 581934 112874 617378
rect 112294 581698 112466 581934
rect 112702 581698 112874 581934
rect 112294 581614 112874 581698
rect 112294 581378 112466 581614
rect 112702 581378 112874 581614
rect 112294 545934 112874 581378
rect 112294 545698 112466 545934
rect 112702 545698 112874 545934
rect 112294 545614 112874 545698
rect 112294 545378 112466 545614
rect 112702 545378 112874 545614
rect 112294 509934 112874 545378
rect 112294 509698 112466 509934
rect 112702 509698 112874 509934
rect 112294 509614 112874 509698
rect 112294 509378 112466 509614
rect 112702 509378 112874 509614
rect 112294 473934 112874 509378
rect 112294 473698 112466 473934
rect 112702 473698 112874 473934
rect 112294 473614 112874 473698
rect 112294 473378 112466 473614
rect 112702 473378 112874 473614
rect 112294 437934 112874 473378
rect 112294 437698 112466 437934
rect 112702 437698 112874 437934
rect 112294 437614 112874 437698
rect 112294 437378 112466 437614
rect 112702 437378 112874 437614
rect 112294 401934 112874 437378
rect 112294 401698 112466 401934
rect 112702 401698 112874 401934
rect 112294 401614 112874 401698
rect 112294 401378 112466 401614
rect 112702 401378 112874 401614
rect 112294 365934 112874 401378
rect 112294 365698 112466 365934
rect 112702 365698 112874 365934
rect 112294 365614 112874 365698
rect 112294 365378 112466 365614
rect 112702 365378 112874 365614
rect 112294 329934 112874 365378
rect 112294 329698 112466 329934
rect 112702 329698 112874 329934
rect 112294 329614 112874 329698
rect 112294 329378 112466 329614
rect 112702 329378 112874 329614
rect 112294 293934 112874 329378
rect 112294 293698 112466 293934
rect 112702 293698 112874 293934
rect 112294 293614 112874 293698
rect 112294 293378 112466 293614
rect 112702 293378 112874 293614
rect 112294 257934 112874 293378
rect 112294 257698 112466 257934
rect 112702 257698 112874 257934
rect 112294 257614 112874 257698
rect 112294 257378 112466 257614
rect 112702 257378 112874 257614
rect 112294 221934 112874 257378
rect 112294 221698 112466 221934
rect 112702 221698 112874 221934
rect 112294 221614 112874 221698
rect 112294 221378 112466 221614
rect 112702 221378 112874 221614
rect 112294 185934 112874 221378
rect 112294 185698 112466 185934
rect 112702 185698 112874 185934
rect 112294 185614 112874 185698
rect 112294 185378 112466 185614
rect 112702 185378 112874 185614
rect 112294 149934 112874 185378
rect 112294 149698 112466 149934
rect 112702 149698 112874 149934
rect 112294 149614 112874 149698
rect 112294 149378 112466 149614
rect 112702 149378 112874 149614
rect 112294 113934 112874 149378
rect 112294 113698 112466 113934
rect 112702 113698 112874 113934
rect 112294 113614 112874 113698
rect 112294 113378 112466 113614
rect 112702 113378 112874 113614
rect 112294 77934 112874 113378
rect 112294 77698 112466 77934
rect 112702 77698 112874 77934
rect 112294 77614 112874 77698
rect 112294 77378 112466 77614
rect 112702 77378 112874 77614
rect 112294 41934 112874 77378
rect 112294 41698 112466 41934
rect 112702 41698 112874 41934
rect 112294 41614 112874 41698
rect 112294 41378 112466 41614
rect 112702 41378 112874 41614
rect 112294 5934 112874 41378
rect 112294 5698 112466 5934
rect 112702 5698 112874 5934
rect 112294 5614 112874 5698
rect 112294 5378 112466 5614
rect 112702 5378 112874 5614
rect 112294 -2186 112874 5378
rect 112294 -2422 112466 -2186
rect 112702 -2422 112874 -2186
rect 112294 -2506 112874 -2422
rect 112294 -2742 112466 -2506
rect 112702 -2742 112874 -2506
rect 112294 -3674 112874 -2742
rect 115774 693414 116354 707962
rect 115774 693178 115946 693414
rect 116182 693178 116354 693414
rect 115774 693094 116354 693178
rect 115774 692858 115946 693094
rect 116182 692858 116354 693094
rect 115774 657414 116354 692858
rect 115774 657178 115946 657414
rect 116182 657178 116354 657414
rect 115774 657094 116354 657178
rect 115774 656858 115946 657094
rect 116182 656858 116354 657094
rect 115774 621414 116354 656858
rect 115774 621178 115946 621414
rect 116182 621178 116354 621414
rect 115774 621094 116354 621178
rect 115774 620858 115946 621094
rect 116182 620858 116354 621094
rect 115774 585414 116354 620858
rect 115774 585178 115946 585414
rect 116182 585178 116354 585414
rect 115774 585094 116354 585178
rect 115774 584858 115946 585094
rect 116182 584858 116354 585094
rect 115774 549414 116354 584858
rect 115774 549178 115946 549414
rect 116182 549178 116354 549414
rect 115774 549094 116354 549178
rect 115774 548858 115946 549094
rect 116182 548858 116354 549094
rect 115774 513414 116354 548858
rect 115774 513178 115946 513414
rect 116182 513178 116354 513414
rect 115774 513094 116354 513178
rect 115774 512858 115946 513094
rect 116182 512858 116354 513094
rect 115774 477414 116354 512858
rect 115774 477178 115946 477414
rect 116182 477178 116354 477414
rect 115774 477094 116354 477178
rect 115774 476858 115946 477094
rect 116182 476858 116354 477094
rect 115774 441414 116354 476858
rect 115774 441178 115946 441414
rect 116182 441178 116354 441414
rect 115774 441094 116354 441178
rect 115774 440858 115946 441094
rect 116182 440858 116354 441094
rect 115774 405414 116354 440858
rect 115774 405178 115946 405414
rect 116182 405178 116354 405414
rect 115774 405094 116354 405178
rect 115774 404858 115946 405094
rect 116182 404858 116354 405094
rect 115774 369414 116354 404858
rect 115774 369178 115946 369414
rect 116182 369178 116354 369414
rect 115774 369094 116354 369178
rect 115774 368858 115946 369094
rect 116182 368858 116354 369094
rect 115774 333414 116354 368858
rect 115774 333178 115946 333414
rect 116182 333178 116354 333414
rect 115774 333094 116354 333178
rect 115774 332858 115946 333094
rect 116182 332858 116354 333094
rect 115774 297414 116354 332858
rect 115774 297178 115946 297414
rect 116182 297178 116354 297414
rect 115774 297094 116354 297178
rect 115774 296858 115946 297094
rect 116182 296858 116354 297094
rect 115774 261414 116354 296858
rect 115774 261178 115946 261414
rect 116182 261178 116354 261414
rect 115774 261094 116354 261178
rect 115774 260858 115946 261094
rect 116182 260858 116354 261094
rect 115774 225414 116354 260858
rect 115774 225178 115946 225414
rect 116182 225178 116354 225414
rect 115774 225094 116354 225178
rect 115774 224858 115946 225094
rect 116182 224858 116354 225094
rect 115774 189414 116354 224858
rect 115774 189178 115946 189414
rect 116182 189178 116354 189414
rect 115774 189094 116354 189178
rect 115774 188858 115946 189094
rect 116182 188858 116354 189094
rect 115774 153414 116354 188858
rect 115774 153178 115946 153414
rect 116182 153178 116354 153414
rect 115774 153094 116354 153178
rect 115774 152858 115946 153094
rect 116182 152858 116354 153094
rect 115774 117414 116354 152858
rect 115774 117178 115946 117414
rect 116182 117178 116354 117414
rect 115774 117094 116354 117178
rect 115774 116858 115946 117094
rect 116182 116858 116354 117094
rect 115774 81414 116354 116858
rect 115774 81178 115946 81414
rect 116182 81178 116354 81414
rect 115774 81094 116354 81178
rect 115774 80858 115946 81094
rect 116182 80858 116354 81094
rect 115774 45414 116354 80858
rect 115774 45178 115946 45414
rect 116182 45178 116354 45414
rect 115774 45094 116354 45178
rect 115774 44858 115946 45094
rect 116182 44858 116354 45094
rect 115774 9414 116354 44858
rect 115774 9178 115946 9414
rect 116182 9178 116354 9414
rect 115774 9094 116354 9178
rect 115774 8858 115946 9094
rect 116182 8858 116354 9094
rect 115774 -4026 116354 8858
rect 115774 -4262 115946 -4026
rect 116182 -4262 116354 -4026
rect 115774 -4346 116354 -4262
rect 115774 -4582 115946 -4346
rect 116182 -4582 116354 -4346
rect 115774 -5514 116354 -4582
rect 119254 696894 119834 709802
rect 137254 711278 137834 711290
rect 137254 711042 137426 711278
rect 137662 711042 137834 711278
rect 137254 710958 137834 711042
rect 137254 710722 137426 710958
rect 137662 710722 137834 710958
rect 133774 709438 134354 709450
rect 133774 709202 133946 709438
rect 134182 709202 134354 709438
rect 133774 709118 134354 709202
rect 133774 708882 133946 709118
rect 134182 708882 134354 709118
rect 130294 707598 130874 707610
rect 130294 707362 130466 707598
rect 130702 707362 130874 707598
rect 130294 707278 130874 707362
rect 130294 707042 130466 707278
rect 130702 707042 130874 707278
rect 119254 696658 119426 696894
rect 119662 696658 119834 696894
rect 119254 696574 119834 696658
rect 119254 696338 119426 696574
rect 119662 696338 119834 696574
rect 119254 660894 119834 696338
rect 119254 660658 119426 660894
rect 119662 660658 119834 660894
rect 119254 660574 119834 660658
rect 119254 660338 119426 660574
rect 119662 660338 119834 660574
rect 119254 624894 119834 660338
rect 119254 624658 119426 624894
rect 119662 624658 119834 624894
rect 119254 624574 119834 624658
rect 119254 624338 119426 624574
rect 119662 624338 119834 624574
rect 119254 588894 119834 624338
rect 119254 588658 119426 588894
rect 119662 588658 119834 588894
rect 119254 588574 119834 588658
rect 119254 588338 119426 588574
rect 119662 588338 119834 588574
rect 119254 552894 119834 588338
rect 119254 552658 119426 552894
rect 119662 552658 119834 552894
rect 119254 552574 119834 552658
rect 119254 552338 119426 552574
rect 119662 552338 119834 552574
rect 119254 516894 119834 552338
rect 119254 516658 119426 516894
rect 119662 516658 119834 516894
rect 119254 516574 119834 516658
rect 119254 516338 119426 516574
rect 119662 516338 119834 516574
rect 119254 480894 119834 516338
rect 119254 480658 119426 480894
rect 119662 480658 119834 480894
rect 119254 480574 119834 480658
rect 119254 480338 119426 480574
rect 119662 480338 119834 480574
rect 119254 444894 119834 480338
rect 119254 444658 119426 444894
rect 119662 444658 119834 444894
rect 119254 444574 119834 444658
rect 119254 444338 119426 444574
rect 119662 444338 119834 444574
rect 119254 408894 119834 444338
rect 119254 408658 119426 408894
rect 119662 408658 119834 408894
rect 119254 408574 119834 408658
rect 119254 408338 119426 408574
rect 119662 408338 119834 408574
rect 119254 372894 119834 408338
rect 119254 372658 119426 372894
rect 119662 372658 119834 372894
rect 119254 372574 119834 372658
rect 119254 372338 119426 372574
rect 119662 372338 119834 372574
rect 119254 336894 119834 372338
rect 119254 336658 119426 336894
rect 119662 336658 119834 336894
rect 119254 336574 119834 336658
rect 119254 336338 119426 336574
rect 119662 336338 119834 336574
rect 119254 300894 119834 336338
rect 119254 300658 119426 300894
rect 119662 300658 119834 300894
rect 119254 300574 119834 300658
rect 119254 300338 119426 300574
rect 119662 300338 119834 300574
rect 119254 264894 119834 300338
rect 119254 264658 119426 264894
rect 119662 264658 119834 264894
rect 119254 264574 119834 264658
rect 119254 264338 119426 264574
rect 119662 264338 119834 264574
rect 119254 228894 119834 264338
rect 119254 228658 119426 228894
rect 119662 228658 119834 228894
rect 119254 228574 119834 228658
rect 119254 228338 119426 228574
rect 119662 228338 119834 228574
rect 119254 192894 119834 228338
rect 119254 192658 119426 192894
rect 119662 192658 119834 192894
rect 119254 192574 119834 192658
rect 119254 192338 119426 192574
rect 119662 192338 119834 192574
rect 119254 156894 119834 192338
rect 119254 156658 119426 156894
rect 119662 156658 119834 156894
rect 119254 156574 119834 156658
rect 119254 156338 119426 156574
rect 119662 156338 119834 156574
rect 119254 120894 119834 156338
rect 119254 120658 119426 120894
rect 119662 120658 119834 120894
rect 119254 120574 119834 120658
rect 119254 120338 119426 120574
rect 119662 120338 119834 120574
rect 119254 84894 119834 120338
rect 119254 84658 119426 84894
rect 119662 84658 119834 84894
rect 119254 84574 119834 84658
rect 119254 84338 119426 84574
rect 119662 84338 119834 84574
rect 119254 48894 119834 84338
rect 119254 48658 119426 48894
rect 119662 48658 119834 48894
rect 119254 48574 119834 48658
rect 119254 48338 119426 48574
rect 119662 48338 119834 48574
rect 119254 12894 119834 48338
rect 119254 12658 119426 12894
rect 119662 12658 119834 12894
rect 119254 12574 119834 12658
rect 119254 12338 119426 12574
rect 119662 12338 119834 12574
rect 101254 -7022 101426 -6786
rect 101662 -7022 101834 -6786
rect 101254 -7106 101834 -7022
rect 101254 -7342 101426 -7106
rect 101662 -7342 101834 -7106
rect 101254 -7354 101834 -7342
rect 119254 -5866 119834 12338
rect 126814 705758 127394 705770
rect 126814 705522 126986 705758
rect 127222 705522 127394 705758
rect 126814 705438 127394 705522
rect 126814 705202 126986 705438
rect 127222 705202 127394 705438
rect 126814 668454 127394 705202
rect 126814 668218 126986 668454
rect 127222 668218 127394 668454
rect 126814 668134 127394 668218
rect 126814 667898 126986 668134
rect 127222 667898 127394 668134
rect 126814 632454 127394 667898
rect 126814 632218 126986 632454
rect 127222 632218 127394 632454
rect 126814 632134 127394 632218
rect 126814 631898 126986 632134
rect 127222 631898 127394 632134
rect 126814 596454 127394 631898
rect 126814 596218 126986 596454
rect 127222 596218 127394 596454
rect 126814 596134 127394 596218
rect 126814 595898 126986 596134
rect 127222 595898 127394 596134
rect 126814 560454 127394 595898
rect 126814 560218 126986 560454
rect 127222 560218 127394 560454
rect 126814 560134 127394 560218
rect 126814 559898 126986 560134
rect 127222 559898 127394 560134
rect 126814 524454 127394 559898
rect 126814 524218 126986 524454
rect 127222 524218 127394 524454
rect 126814 524134 127394 524218
rect 126814 523898 126986 524134
rect 127222 523898 127394 524134
rect 126814 488454 127394 523898
rect 126814 488218 126986 488454
rect 127222 488218 127394 488454
rect 126814 488134 127394 488218
rect 126814 487898 126986 488134
rect 127222 487898 127394 488134
rect 126814 452454 127394 487898
rect 126814 452218 126986 452454
rect 127222 452218 127394 452454
rect 126814 452134 127394 452218
rect 126814 451898 126986 452134
rect 127222 451898 127394 452134
rect 126814 416454 127394 451898
rect 126814 416218 126986 416454
rect 127222 416218 127394 416454
rect 126814 416134 127394 416218
rect 126814 415898 126986 416134
rect 127222 415898 127394 416134
rect 126814 380454 127394 415898
rect 126814 380218 126986 380454
rect 127222 380218 127394 380454
rect 126814 380134 127394 380218
rect 126814 379898 126986 380134
rect 127222 379898 127394 380134
rect 126814 344454 127394 379898
rect 126814 344218 126986 344454
rect 127222 344218 127394 344454
rect 126814 344134 127394 344218
rect 126814 343898 126986 344134
rect 127222 343898 127394 344134
rect 126814 308454 127394 343898
rect 126814 308218 126986 308454
rect 127222 308218 127394 308454
rect 126814 308134 127394 308218
rect 126814 307898 126986 308134
rect 127222 307898 127394 308134
rect 126814 272454 127394 307898
rect 126814 272218 126986 272454
rect 127222 272218 127394 272454
rect 126814 272134 127394 272218
rect 126814 271898 126986 272134
rect 127222 271898 127394 272134
rect 126814 236454 127394 271898
rect 126814 236218 126986 236454
rect 127222 236218 127394 236454
rect 126814 236134 127394 236218
rect 126814 235898 126986 236134
rect 127222 235898 127394 236134
rect 126814 200454 127394 235898
rect 126814 200218 126986 200454
rect 127222 200218 127394 200454
rect 126814 200134 127394 200218
rect 126814 199898 126986 200134
rect 127222 199898 127394 200134
rect 126814 164454 127394 199898
rect 126814 164218 126986 164454
rect 127222 164218 127394 164454
rect 126814 164134 127394 164218
rect 126814 163898 126986 164134
rect 127222 163898 127394 164134
rect 126814 128454 127394 163898
rect 126814 128218 126986 128454
rect 127222 128218 127394 128454
rect 126814 128134 127394 128218
rect 126814 127898 126986 128134
rect 127222 127898 127394 128134
rect 126814 92454 127394 127898
rect 126814 92218 126986 92454
rect 127222 92218 127394 92454
rect 126814 92134 127394 92218
rect 126814 91898 126986 92134
rect 127222 91898 127394 92134
rect 126814 56454 127394 91898
rect 126814 56218 126986 56454
rect 127222 56218 127394 56454
rect 126814 56134 127394 56218
rect 126814 55898 126986 56134
rect 127222 55898 127394 56134
rect 126814 20454 127394 55898
rect 126814 20218 126986 20454
rect 127222 20218 127394 20454
rect 126814 20134 127394 20218
rect 126814 19898 126986 20134
rect 127222 19898 127394 20134
rect 126814 -1266 127394 19898
rect 126814 -1502 126986 -1266
rect 127222 -1502 127394 -1266
rect 126814 -1586 127394 -1502
rect 126814 -1822 126986 -1586
rect 127222 -1822 127394 -1586
rect 126814 -1834 127394 -1822
rect 130294 671934 130874 707042
rect 130294 671698 130466 671934
rect 130702 671698 130874 671934
rect 130294 671614 130874 671698
rect 130294 671378 130466 671614
rect 130702 671378 130874 671614
rect 130294 635934 130874 671378
rect 130294 635698 130466 635934
rect 130702 635698 130874 635934
rect 130294 635614 130874 635698
rect 130294 635378 130466 635614
rect 130702 635378 130874 635614
rect 130294 599934 130874 635378
rect 130294 599698 130466 599934
rect 130702 599698 130874 599934
rect 130294 599614 130874 599698
rect 130294 599378 130466 599614
rect 130702 599378 130874 599614
rect 130294 563934 130874 599378
rect 130294 563698 130466 563934
rect 130702 563698 130874 563934
rect 130294 563614 130874 563698
rect 130294 563378 130466 563614
rect 130702 563378 130874 563614
rect 130294 527934 130874 563378
rect 130294 527698 130466 527934
rect 130702 527698 130874 527934
rect 130294 527614 130874 527698
rect 130294 527378 130466 527614
rect 130702 527378 130874 527614
rect 130294 491934 130874 527378
rect 130294 491698 130466 491934
rect 130702 491698 130874 491934
rect 130294 491614 130874 491698
rect 130294 491378 130466 491614
rect 130702 491378 130874 491614
rect 130294 455934 130874 491378
rect 130294 455698 130466 455934
rect 130702 455698 130874 455934
rect 130294 455614 130874 455698
rect 130294 455378 130466 455614
rect 130702 455378 130874 455614
rect 130294 419934 130874 455378
rect 130294 419698 130466 419934
rect 130702 419698 130874 419934
rect 130294 419614 130874 419698
rect 130294 419378 130466 419614
rect 130702 419378 130874 419614
rect 130294 383934 130874 419378
rect 130294 383698 130466 383934
rect 130702 383698 130874 383934
rect 130294 383614 130874 383698
rect 130294 383378 130466 383614
rect 130702 383378 130874 383614
rect 130294 347934 130874 383378
rect 130294 347698 130466 347934
rect 130702 347698 130874 347934
rect 130294 347614 130874 347698
rect 130294 347378 130466 347614
rect 130702 347378 130874 347614
rect 130294 311934 130874 347378
rect 130294 311698 130466 311934
rect 130702 311698 130874 311934
rect 130294 311614 130874 311698
rect 130294 311378 130466 311614
rect 130702 311378 130874 311614
rect 130294 275934 130874 311378
rect 130294 275698 130466 275934
rect 130702 275698 130874 275934
rect 130294 275614 130874 275698
rect 130294 275378 130466 275614
rect 130702 275378 130874 275614
rect 130294 239934 130874 275378
rect 130294 239698 130466 239934
rect 130702 239698 130874 239934
rect 130294 239614 130874 239698
rect 130294 239378 130466 239614
rect 130702 239378 130874 239614
rect 130294 203934 130874 239378
rect 130294 203698 130466 203934
rect 130702 203698 130874 203934
rect 130294 203614 130874 203698
rect 130294 203378 130466 203614
rect 130702 203378 130874 203614
rect 130294 167934 130874 203378
rect 130294 167698 130466 167934
rect 130702 167698 130874 167934
rect 130294 167614 130874 167698
rect 130294 167378 130466 167614
rect 130702 167378 130874 167614
rect 130294 131934 130874 167378
rect 130294 131698 130466 131934
rect 130702 131698 130874 131934
rect 130294 131614 130874 131698
rect 130294 131378 130466 131614
rect 130702 131378 130874 131614
rect 130294 95934 130874 131378
rect 130294 95698 130466 95934
rect 130702 95698 130874 95934
rect 130294 95614 130874 95698
rect 130294 95378 130466 95614
rect 130702 95378 130874 95614
rect 130294 59934 130874 95378
rect 130294 59698 130466 59934
rect 130702 59698 130874 59934
rect 130294 59614 130874 59698
rect 130294 59378 130466 59614
rect 130702 59378 130874 59614
rect 130294 23934 130874 59378
rect 130294 23698 130466 23934
rect 130702 23698 130874 23934
rect 130294 23614 130874 23698
rect 130294 23378 130466 23614
rect 130702 23378 130874 23614
rect 130294 -3106 130874 23378
rect 130294 -3342 130466 -3106
rect 130702 -3342 130874 -3106
rect 130294 -3426 130874 -3342
rect 130294 -3662 130466 -3426
rect 130702 -3662 130874 -3426
rect 130294 -3674 130874 -3662
rect 133774 675414 134354 708882
rect 133774 675178 133946 675414
rect 134182 675178 134354 675414
rect 133774 675094 134354 675178
rect 133774 674858 133946 675094
rect 134182 674858 134354 675094
rect 133774 639414 134354 674858
rect 133774 639178 133946 639414
rect 134182 639178 134354 639414
rect 133774 639094 134354 639178
rect 133774 638858 133946 639094
rect 134182 638858 134354 639094
rect 133774 603414 134354 638858
rect 133774 603178 133946 603414
rect 134182 603178 134354 603414
rect 133774 603094 134354 603178
rect 133774 602858 133946 603094
rect 134182 602858 134354 603094
rect 133774 567414 134354 602858
rect 133774 567178 133946 567414
rect 134182 567178 134354 567414
rect 133774 567094 134354 567178
rect 133774 566858 133946 567094
rect 134182 566858 134354 567094
rect 133774 531414 134354 566858
rect 133774 531178 133946 531414
rect 134182 531178 134354 531414
rect 133774 531094 134354 531178
rect 133774 530858 133946 531094
rect 134182 530858 134354 531094
rect 133774 495414 134354 530858
rect 133774 495178 133946 495414
rect 134182 495178 134354 495414
rect 133774 495094 134354 495178
rect 133774 494858 133946 495094
rect 134182 494858 134354 495094
rect 133774 459414 134354 494858
rect 133774 459178 133946 459414
rect 134182 459178 134354 459414
rect 133774 459094 134354 459178
rect 133774 458858 133946 459094
rect 134182 458858 134354 459094
rect 133774 423414 134354 458858
rect 133774 423178 133946 423414
rect 134182 423178 134354 423414
rect 133774 423094 134354 423178
rect 133774 422858 133946 423094
rect 134182 422858 134354 423094
rect 133774 387414 134354 422858
rect 133774 387178 133946 387414
rect 134182 387178 134354 387414
rect 133774 387094 134354 387178
rect 133774 386858 133946 387094
rect 134182 386858 134354 387094
rect 133774 351414 134354 386858
rect 133774 351178 133946 351414
rect 134182 351178 134354 351414
rect 133774 351094 134354 351178
rect 133774 350858 133946 351094
rect 134182 350858 134354 351094
rect 133774 315414 134354 350858
rect 133774 315178 133946 315414
rect 134182 315178 134354 315414
rect 133774 315094 134354 315178
rect 133774 314858 133946 315094
rect 134182 314858 134354 315094
rect 133774 279414 134354 314858
rect 133774 279178 133946 279414
rect 134182 279178 134354 279414
rect 133774 279094 134354 279178
rect 133774 278858 133946 279094
rect 134182 278858 134354 279094
rect 133774 243414 134354 278858
rect 133774 243178 133946 243414
rect 134182 243178 134354 243414
rect 133774 243094 134354 243178
rect 133774 242858 133946 243094
rect 134182 242858 134354 243094
rect 133774 207414 134354 242858
rect 133774 207178 133946 207414
rect 134182 207178 134354 207414
rect 133774 207094 134354 207178
rect 133774 206858 133946 207094
rect 134182 206858 134354 207094
rect 133774 171414 134354 206858
rect 133774 171178 133946 171414
rect 134182 171178 134354 171414
rect 133774 171094 134354 171178
rect 133774 170858 133946 171094
rect 134182 170858 134354 171094
rect 133774 135414 134354 170858
rect 133774 135178 133946 135414
rect 134182 135178 134354 135414
rect 133774 135094 134354 135178
rect 133774 134858 133946 135094
rect 134182 134858 134354 135094
rect 133774 99414 134354 134858
rect 133774 99178 133946 99414
rect 134182 99178 134354 99414
rect 133774 99094 134354 99178
rect 133774 98858 133946 99094
rect 134182 98858 134354 99094
rect 133774 63414 134354 98858
rect 133774 63178 133946 63414
rect 134182 63178 134354 63414
rect 133774 63094 134354 63178
rect 133774 62858 133946 63094
rect 134182 62858 134354 63094
rect 133774 27414 134354 62858
rect 133774 27178 133946 27414
rect 134182 27178 134354 27414
rect 133774 27094 134354 27178
rect 133774 26858 133946 27094
rect 134182 26858 134354 27094
rect 133774 -4946 134354 26858
rect 133774 -5182 133946 -4946
rect 134182 -5182 134354 -4946
rect 133774 -5266 134354 -5182
rect 133774 -5502 133946 -5266
rect 134182 -5502 134354 -5266
rect 133774 -5514 134354 -5502
rect 137254 678894 137834 710722
rect 155254 710358 155834 711290
rect 155254 710122 155426 710358
rect 155662 710122 155834 710358
rect 155254 710038 155834 710122
rect 155254 709802 155426 710038
rect 155662 709802 155834 710038
rect 151774 708518 152354 709450
rect 151774 708282 151946 708518
rect 152182 708282 152354 708518
rect 151774 708198 152354 708282
rect 151774 707962 151946 708198
rect 152182 707962 152354 708198
rect 148294 706678 148874 707610
rect 148294 706442 148466 706678
rect 148702 706442 148874 706678
rect 148294 706358 148874 706442
rect 148294 706122 148466 706358
rect 148702 706122 148874 706358
rect 137254 678658 137426 678894
rect 137662 678658 137834 678894
rect 137254 678574 137834 678658
rect 137254 678338 137426 678574
rect 137662 678338 137834 678574
rect 137254 642894 137834 678338
rect 137254 642658 137426 642894
rect 137662 642658 137834 642894
rect 137254 642574 137834 642658
rect 137254 642338 137426 642574
rect 137662 642338 137834 642574
rect 137254 606894 137834 642338
rect 137254 606658 137426 606894
rect 137662 606658 137834 606894
rect 137254 606574 137834 606658
rect 137254 606338 137426 606574
rect 137662 606338 137834 606574
rect 137254 570894 137834 606338
rect 137254 570658 137426 570894
rect 137662 570658 137834 570894
rect 137254 570574 137834 570658
rect 137254 570338 137426 570574
rect 137662 570338 137834 570574
rect 137254 534894 137834 570338
rect 137254 534658 137426 534894
rect 137662 534658 137834 534894
rect 137254 534574 137834 534658
rect 137254 534338 137426 534574
rect 137662 534338 137834 534574
rect 137254 498894 137834 534338
rect 137254 498658 137426 498894
rect 137662 498658 137834 498894
rect 137254 498574 137834 498658
rect 137254 498338 137426 498574
rect 137662 498338 137834 498574
rect 137254 462894 137834 498338
rect 137254 462658 137426 462894
rect 137662 462658 137834 462894
rect 137254 462574 137834 462658
rect 137254 462338 137426 462574
rect 137662 462338 137834 462574
rect 137254 426894 137834 462338
rect 137254 426658 137426 426894
rect 137662 426658 137834 426894
rect 137254 426574 137834 426658
rect 137254 426338 137426 426574
rect 137662 426338 137834 426574
rect 137254 390894 137834 426338
rect 137254 390658 137426 390894
rect 137662 390658 137834 390894
rect 137254 390574 137834 390658
rect 137254 390338 137426 390574
rect 137662 390338 137834 390574
rect 137254 354894 137834 390338
rect 137254 354658 137426 354894
rect 137662 354658 137834 354894
rect 137254 354574 137834 354658
rect 137254 354338 137426 354574
rect 137662 354338 137834 354574
rect 137254 318894 137834 354338
rect 137254 318658 137426 318894
rect 137662 318658 137834 318894
rect 137254 318574 137834 318658
rect 137254 318338 137426 318574
rect 137662 318338 137834 318574
rect 137254 282894 137834 318338
rect 137254 282658 137426 282894
rect 137662 282658 137834 282894
rect 137254 282574 137834 282658
rect 137254 282338 137426 282574
rect 137662 282338 137834 282574
rect 137254 246894 137834 282338
rect 137254 246658 137426 246894
rect 137662 246658 137834 246894
rect 137254 246574 137834 246658
rect 137254 246338 137426 246574
rect 137662 246338 137834 246574
rect 137254 210894 137834 246338
rect 137254 210658 137426 210894
rect 137662 210658 137834 210894
rect 137254 210574 137834 210658
rect 137254 210338 137426 210574
rect 137662 210338 137834 210574
rect 137254 174894 137834 210338
rect 137254 174658 137426 174894
rect 137662 174658 137834 174894
rect 137254 174574 137834 174658
rect 137254 174338 137426 174574
rect 137662 174338 137834 174574
rect 137254 138894 137834 174338
rect 137254 138658 137426 138894
rect 137662 138658 137834 138894
rect 137254 138574 137834 138658
rect 137254 138338 137426 138574
rect 137662 138338 137834 138574
rect 137254 102894 137834 138338
rect 137254 102658 137426 102894
rect 137662 102658 137834 102894
rect 137254 102574 137834 102658
rect 137254 102338 137426 102574
rect 137662 102338 137834 102574
rect 137254 66894 137834 102338
rect 137254 66658 137426 66894
rect 137662 66658 137834 66894
rect 137254 66574 137834 66658
rect 137254 66338 137426 66574
rect 137662 66338 137834 66574
rect 137254 30894 137834 66338
rect 137254 30658 137426 30894
rect 137662 30658 137834 30894
rect 137254 30574 137834 30658
rect 137254 30338 137426 30574
rect 137662 30338 137834 30574
rect 119254 -6102 119426 -5866
rect 119662 -6102 119834 -5866
rect 119254 -6186 119834 -6102
rect 119254 -6422 119426 -6186
rect 119662 -6422 119834 -6186
rect 119254 -7354 119834 -6422
rect 137254 -6786 137834 30338
rect 144814 704838 145394 705770
rect 144814 704602 144986 704838
rect 145222 704602 145394 704838
rect 144814 704518 145394 704602
rect 144814 704282 144986 704518
rect 145222 704282 145394 704518
rect 144814 686454 145394 704282
rect 144814 686218 144986 686454
rect 145222 686218 145394 686454
rect 144814 686134 145394 686218
rect 144814 685898 144986 686134
rect 145222 685898 145394 686134
rect 144814 650454 145394 685898
rect 144814 650218 144986 650454
rect 145222 650218 145394 650454
rect 144814 650134 145394 650218
rect 144814 649898 144986 650134
rect 145222 649898 145394 650134
rect 144814 614454 145394 649898
rect 144814 614218 144986 614454
rect 145222 614218 145394 614454
rect 144814 614134 145394 614218
rect 144814 613898 144986 614134
rect 145222 613898 145394 614134
rect 144814 578454 145394 613898
rect 144814 578218 144986 578454
rect 145222 578218 145394 578454
rect 144814 578134 145394 578218
rect 144814 577898 144986 578134
rect 145222 577898 145394 578134
rect 144814 542454 145394 577898
rect 144814 542218 144986 542454
rect 145222 542218 145394 542454
rect 144814 542134 145394 542218
rect 144814 541898 144986 542134
rect 145222 541898 145394 542134
rect 144814 506454 145394 541898
rect 144814 506218 144986 506454
rect 145222 506218 145394 506454
rect 144814 506134 145394 506218
rect 144814 505898 144986 506134
rect 145222 505898 145394 506134
rect 144814 470454 145394 505898
rect 144814 470218 144986 470454
rect 145222 470218 145394 470454
rect 144814 470134 145394 470218
rect 144814 469898 144986 470134
rect 145222 469898 145394 470134
rect 144814 434454 145394 469898
rect 144814 434218 144986 434454
rect 145222 434218 145394 434454
rect 144814 434134 145394 434218
rect 144814 433898 144986 434134
rect 145222 433898 145394 434134
rect 144814 398454 145394 433898
rect 144814 398218 144986 398454
rect 145222 398218 145394 398454
rect 144814 398134 145394 398218
rect 144814 397898 144986 398134
rect 145222 397898 145394 398134
rect 144814 362454 145394 397898
rect 144814 362218 144986 362454
rect 145222 362218 145394 362454
rect 144814 362134 145394 362218
rect 144814 361898 144986 362134
rect 145222 361898 145394 362134
rect 144814 326454 145394 361898
rect 144814 326218 144986 326454
rect 145222 326218 145394 326454
rect 144814 326134 145394 326218
rect 144814 325898 144986 326134
rect 145222 325898 145394 326134
rect 144814 290454 145394 325898
rect 144814 290218 144986 290454
rect 145222 290218 145394 290454
rect 144814 290134 145394 290218
rect 144814 289898 144986 290134
rect 145222 289898 145394 290134
rect 144814 254454 145394 289898
rect 144814 254218 144986 254454
rect 145222 254218 145394 254454
rect 144814 254134 145394 254218
rect 144814 253898 144986 254134
rect 145222 253898 145394 254134
rect 144814 218454 145394 253898
rect 144814 218218 144986 218454
rect 145222 218218 145394 218454
rect 144814 218134 145394 218218
rect 144814 217898 144986 218134
rect 145222 217898 145394 218134
rect 144814 182454 145394 217898
rect 144814 182218 144986 182454
rect 145222 182218 145394 182454
rect 144814 182134 145394 182218
rect 144814 181898 144986 182134
rect 145222 181898 145394 182134
rect 144814 146454 145394 181898
rect 144814 146218 144986 146454
rect 145222 146218 145394 146454
rect 144814 146134 145394 146218
rect 144814 145898 144986 146134
rect 145222 145898 145394 146134
rect 144814 110454 145394 145898
rect 144814 110218 144986 110454
rect 145222 110218 145394 110454
rect 144814 110134 145394 110218
rect 144814 109898 144986 110134
rect 145222 109898 145394 110134
rect 144814 74454 145394 109898
rect 144814 74218 144986 74454
rect 145222 74218 145394 74454
rect 144814 74134 145394 74218
rect 144814 73898 144986 74134
rect 145222 73898 145394 74134
rect 144814 38454 145394 73898
rect 144814 38218 144986 38454
rect 145222 38218 145394 38454
rect 144814 38134 145394 38218
rect 144814 37898 144986 38134
rect 145222 37898 145394 38134
rect 144814 2454 145394 37898
rect 144814 2218 144986 2454
rect 145222 2218 145394 2454
rect 144814 2134 145394 2218
rect 144814 1898 144986 2134
rect 145222 1898 145394 2134
rect 144814 -346 145394 1898
rect 144814 -582 144986 -346
rect 145222 -582 145394 -346
rect 144814 -666 145394 -582
rect 144814 -902 144986 -666
rect 145222 -902 145394 -666
rect 144814 -1834 145394 -902
rect 148294 689934 148874 706122
rect 148294 689698 148466 689934
rect 148702 689698 148874 689934
rect 148294 689614 148874 689698
rect 148294 689378 148466 689614
rect 148702 689378 148874 689614
rect 148294 653934 148874 689378
rect 148294 653698 148466 653934
rect 148702 653698 148874 653934
rect 148294 653614 148874 653698
rect 148294 653378 148466 653614
rect 148702 653378 148874 653614
rect 148294 617934 148874 653378
rect 148294 617698 148466 617934
rect 148702 617698 148874 617934
rect 148294 617614 148874 617698
rect 148294 617378 148466 617614
rect 148702 617378 148874 617614
rect 148294 581934 148874 617378
rect 148294 581698 148466 581934
rect 148702 581698 148874 581934
rect 148294 581614 148874 581698
rect 148294 581378 148466 581614
rect 148702 581378 148874 581614
rect 148294 545934 148874 581378
rect 148294 545698 148466 545934
rect 148702 545698 148874 545934
rect 148294 545614 148874 545698
rect 148294 545378 148466 545614
rect 148702 545378 148874 545614
rect 148294 509934 148874 545378
rect 148294 509698 148466 509934
rect 148702 509698 148874 509934
rect 148294 509614 148874 509698
rect 148294 509378 148466 509614
rect 148702 509378 148874 509614
rect 148294 473934 148874 509378
rect 148294 473698 148466 473934
rect 148702 473698 148874 473934
rect 148294 473614 148874 473698
rect 148294 473378 148466 473614
rect 148702 473378 148874 473614
rect 148294 437934 148874 473378
rect 148294 437698 148466 437934
rect 148702 437698 148874 437934
rect 148294 437614 148874 437698
rect 148294 437378 148466 437614
rect 148702 437378 148874 437614
rect 148294 401934 148874 437378
rect 148294 401698 148466 401934
rect 148702 401698 148874 401934
rect 148294 401614 148874 401698
rect 148294 401378 148466 401614
rect 148702 401378 148874 401614
rect 148294 365934 148874 401378
rect 148294 365698 148466 365934
rect 148702 365698 148874 365934
rect 148294 365614 148874 365698
rect 148294 365378 148466 365614
rect 148702 365378 148874 365614
rect 148294 329934 148874 365378
rect 148294 329698 148466 329934
rect 148702 329698 148874 329934
rect 148294 329614 148874 329698
rect 148294 329378 148466 329614
rect 148702 329378 148874 329614
rect 148294 293934 148874 329378
rect 148294 293698 148466 293934
rect 148702 293698 148874 293934
rect 148294 293614 148874 293698
rect 148294 293378 148466 293614
rect 148702 293378 148874 293614
rect 148294 257934 148874 293378
rect 148294 257698 148466 257934
rect 148702 257698 148874 257934
rect 148294 257614 148874 257698
rect 148294 257378 148466 257614
rect 148702 257378 148874 257614
rect 148294 221934 148874 257378
rect 148294 221698 148466 221934
rect 148702 221698 148874 221934
rect 148294 221614 148874 221698
rect 148294 221378 148466 221614
rect 148702 221378 148874 221614
rect 148294 185934 148874 221378
rect 148294 185698 148466 185934
rect 148702 185698 148874 185934
rect 148294 185614 148874 185698
rect 148294 185378 148466 185614
rect 148702 185378 148874 185614
rect 148294 149934 148874 185378
rect 148294 149698 148466 149934
rect 148702 149698 148874 149934
rect 148294 149614 148874 149698
rect 148294 149378 148466 149614
rect 148702 149378 148874 149614
rect 148294 113934 148874 149378
rect 148294 113698 148466 113934
rect 148702 113698 148874 113934
rect 148294 113614 148874 113698
rect 148294 113378 148466 113614
rect 148702 113378 148874 113614
rect 148294 77934 148874 113378
rect 148294 77698 148466 77934
rect 148702 77698 148874 77934
rect 148294 77614 148874 77698
rect 148294 77378 148466 77614
rect 148702 77378 148874 77614
rect 148294 41934 148874 77378
rect 148294 41698 148466 41934
rect 148702 41698 148874 41934
rect 148294 41614 148874 41698
rect 148294 41378 148466 41614
rect 148702 41378 148874 41614
rect 148294 5934 148874 41378
rect 148294 5698 148466 5934
rect 148702 5698 148874 5934
rect 148294 5614 148874 5698
rect 148294 5378 148466 5614
rect 148702 5378 148874 5614
rect 148294 -2186 148874 5378
rect 148294 -2422 148466 -2186
rect 148702 -2422 148874 -2186
rect 148294 -2506 148874 -2422
rect 148294 -2742 148466 -2506
rect 148702 -2742 148874 -2506
rect 148294 -3674 148874 -2742
rect 151774 693414 152354 707962
rect 151774 693178 151946 693414
rect 152182 693178 152354 693414
rect 151774 693094 152354 693178
rect 151774 692858 151946 693094
rect 152182 692858 152354 693094
rect 151774 657414 152354 692858
rect 151774 657178 151946 657414
rect 152182 657178 152354 657414
rect 151774 657094 152354 657178
rect 151774 656858 151946 657094
rect 152182 656858 152354 657094
rect 151774 621414 152354 656858
rect 151774 621178 151946 621414
rect 152182 621178 152354 621414
rect 151774 621094 152354 621178
rect 151774 620858 151946 621094
rect 152182 620858 152354 621094
rect 151774 585414 152354 620858
rect 151774 585178 151946 585414
rect 152182 585178 152354 585414
rect 151774 585094 152354 585178
rect 151774 584858 151946 585094
rect 152182 584858 152354 585094
rect 151774 549414 152354 584858
rect 151774 549178 151946 549414
rect 152182 549178 152354 549414
rect 151774 549094 152354 549178
rect 151774 548858 151946 549094
rect 152182 548858 152354 549094
rect 151774 513414 152354 548858
rect 151774 513178 151946 513414
rect 152182 513178 152354 513414
rect 151774 513094 152354 513178
rect 151774 512858 151946 513094
rect 152182 512858 152354 513094
rect 151774 477414 152354 512858
rect 151774 477178 151946 477414
rect 152182 477178 152354 477414
rect 151774 477094 152354 477178
rect 151774 476858 151946 477094
rect 152182 476858 152354 477094
rect 151774 441414 152354 476858
rect 151774 441178 151946 441414
rect 152182 441178 152354 441414
rect 151774 441094 152354 441178
rect 151774 440858 151946 441094
rect 152182 440858 152354 441094
rect 151774 405414 152354 440858
rect 151774 405178 151946 405414
rect 152182 405178 152354 405414
rect 151774 405094 152354 405178
rect 151774 404858 151946 405094
rect 152182 404858 152354 405094
rect 151774 369414 152354 404858
rect 151774 369178 151946 369414
rect 152182 369178 152354 369414
rect 151774 369094 152354 369178
rect 151774 368858 151946 369094
rect 152182 368858 152354 369094
rect 151774 333414 152354 368858
rect 151774 333178 151946 333414
rect 152182 333178 152354 333414
rect 151774 333094 152354 333178
rect 151774 332858 151946 333094
rect 152182 332858 152354 333094
rect 151774 297414 152354 332858
rect 151774 297178 151946 297414
rect 152182 297178 152354 297414
rect 151774 297094 152354 297178
rect 151774 296858 151946 297094
rect 152182 296858 152354 297094
rect 151774 261414 152354 296858
rect 151774 261178 151946 261414
rect 152182 261178 152354 261414
rect 151774 261094 152354 261178
rect 151774 260858 151946 261094
rect 152182 260858 152354 261094
rect 151774 225414 152354 260858
rect 151774 225178 151946 225414
rect 152182 225178 152354 225414
rect 151774 225094 152354 225178
rect 151774 224858 151946 225094
rect 152182 224858 152354 225094
rect 151774 189414 152354 224858
rect 151774 189178 151946 189414
rect 152182 189178 152354 189414
rect 151774 189094 152354 189178
rect 151774 188858 151946 189094
rect 152182 188858 152354 189094
rect 151774 153414 152354 188858
rect 151774 153178 151946 153414
rect 152182 153178 152354 153414
rect 151774 153094 152354 153178
rect 151774 152858 151946 153094
rect 152182 152858 152354 153094
rect 151774 117414 152354 152858
rect 151774 117178 151946 117414
rect 152182 117178 152354 117414
rect 151774 117094 152354 117178
rect 151774 116858 151946 117094
rect 152182 116858 152354 117094
rect 151774 81414 152354 116858
rect 151774 81178 151946 81414
rect 152182 81178 152354 81414
rect 151774 81094 152354 81178
rect 151774 80858 151946 81094
rect 152182 80858 152354 81094
rect 151774 45414 152354 80858
rect 151774 45178 151946 45414
rect 152182 45178 152354 45414
rect 151774 45094 152354 45178
rect 151774 44858 151946 45094
rect 152182 44858 152354 45094
rect 151774 9414 152354 44858
rect 151774 9178 151946 9414
rect 152182 9178 152354 9414
rect 151774 9094 152354 9178
rect 151774 8858 151946 9094
rect 152182 8858 152354 9094
rect 151774 -4026 152354 8858
rect 151774 -4262 151946 -4026
rect 152182 -4262 152354 -4026
rect 151774 -4346 152354 -4262
rect 151774 -4582 151946 -4346
rect 152182 -4582 152354 -4346
rect 151774 -5514 152354 -4582
rect 155254 696894 155834 709802
rect 173254 711278 173834 711290
rect 173254 711042 173426 711278
rect 173662 711042 173834 711278
rect 173254 710958 173834 711042
rect 173254 710722 173426 710958
rect 173662 710722 173834 710958
rect 169774 709438 170354 709450
rect 169774 709202 169946 709438
rect 170182 709202 170354 709438
rect 169774 709118 170354 709202
rect 169774 708882 169946 709118
rect 170182 708882 170354 709118
rect 166294 707598 166874 707610
rect 166294 707362 166466 707598
rect 166702 707362 166874 707598
rect 166294 707278 166874 707362
rect 166294 707042 166466 707278
rect 166702 707042 166874 707278
rect 155254 696658 155426 696894
rect 155662 696658 155834 696894
rect 155254 696574 155834 696658
rect 155254 696338 155426 696574
rect 155662 696338 155834 696574
rect 155254 660894 155834 696338
rect 155254 660658 155426 660894
rect 155662 660658 155834 660894
rect 155254 660574 155834 660658
rect 155254 660338 155426 660574
rect 155662 660338 155834 660574
rect 155254 624894 155834 660338
rect 155254 624658 155426 624894
rect 155662 624658 155834 624894
rect 155254 624574 155834 624658
rect 155254 624338 155426 624574
rect 155662 624338 155834 624574
rect 155254 588894 155834 624338
rect 155254 588658 155426 588894
rect 155662 588658 155834 588894
rect 155254 588574 155834 588658
rect 155254 588338 155426 588574
rect 155662 588338 155834 588574
rect 155254 552894 155834 588338
rect 155254 552658 155426 552894
rect 155662 552658 155834 552894
rect 155254 552574 155834 552658
rect 155254 552338 155426 552574
rect 155662 552338 155834 552574
rect 155254 516894 155834 552338
rect 155254 516658 155426 516894
rect 155662 516658 155834 516894
rect 155254 516574 155834 516658
rect 155254 516338 155426 516574
rect 155662 516338 155834 516574
rect 155254 480894 155834 516338
rect 155254 480658 155426 480894
rect 155662 480658 155834 480894
rect 155254 480574 155834 480658
rect 155254 480338 155426 480574
rect 155662 480338 155834 480574
rect 155254 444894 155834 480338
rect 155254 444658 155426 444894
rect 155662 444658 155834 444894
rect 155254 444574 155834 444658
rect 155254 444338 155426 444574
rect 155662 444338 155834 444574
rect 155254 408894 155834 444338
rect 155254 408658 155426 408894
rect 155662 408658 155834 408894
rect 155254 408574 155834 408658
rect 155254 408338 155426 408574
rect 155662 408338 155834 408574
rect 155254 372894 155834 408338
rect 155254 372658 155426 372894
rect 155662 372658 155834 372894
rect 155254 372574 155834 372658
rect 155254 372338 155426 372574
rect 155662 372338 155834 372574
rect 155254 336894 155834 372338
rect 155254 336658 155426 336894
rect 155662 336658 155834 336894
rect 155254 336574 155834 336658
rect 155254 336338 155426 336574
rect 155662 336338 155834 336574
rect 155254 300894 155834 336338
rect 155254 300658 155426 300894
rect 155662 300658 155834 300894
rect 155254 300574 155834 300658
rect 155254 300338 155426 300574
rect 155662 300338 155834 300574
rect 155254 264894 155834 300338
rect 155254 264658 155426 264894
rect 155662 264658 155834 264894
rect 155254 264574 155834 264658
rect 155254 264338 155426 264574
rect 155662 264338 155834 264574
rect 155254 228894 155834 264338
rect 155254 228658 155426 228894
rect 155662 228658 155834 228894
rect 155254 228574 155834 228658
rect 155254 228338 155426 228574
rect 155662 228338 155834 228574
rect 155254 192894 155834 228338
rect 155254 192658 155426 192894
rect 155662 192658 155834 192894
rect 155254 192574 155834 192658
rect 155254 192338 155426 192574
rect 155662 192338 155834 192574
rect 155254 156894 155834 192338
rect 155254 156658 155426 156894
rect 155662 156658 155834 156894
rect 155254 156574 155834 156658
rect 155254 156338 155426 156574
rect 155662 156338 155834 156574
rect 155254 120894 155834 156338
rect 155254 120658 155426 120894
rect 155662 120658 155834 120894
rect 155254 120574 155834 120658
rect 155254 120338 155426 120574
rect 155662 120338 155834 120574
rect 155254 84894 155834 120338
rect 155254 84658 155426 84894
rect 155662 84658 155834 84894
rect 155254 84574 155834 84658
rect 155254 84338 155426 84574
rect 155662 84338 155834 84574
rect 155254 48894 155834 84338
rect 155254 48658 155426 48894
rect 155662 48658 155834 48894
rect 155254 48574 155834 48658
rect 155254 48338 155426 48574
rect 155662 48338 155834 48574
rect 155254 12894 155834 48338
rect 155254 12658 155426 12894
rect 155662 12658 155834 12894
rect 155254 12574 155834 12658
rect 155254 12338 155426 12574
rect 155662 12338 155834 12574
rect 137254 -7022 137426 -6786
rect 137662 -7022 137834 -6786
rect 137254 -7106 137834 -7022
rect 137254 -7342 137426 -7106
rect 137662 -7342 137834 -7106
rect 137254 -7354 137834 -7342
rect 155254 -5866 155834 12338
rect 162814 705758 163394 705770
rect 162814 705522 162986 705758
rect 163222 705522 163394 705758
rect 162814 705438 163394 705522
rect 162814 705202 162986 705438
rect 163222 705202 163394 705438
rect 162814 668454 163394 705202
rect 162814 668218 162986 668454
rect 163222 668218 163394 668454
rect 162814 668134 163394 668218
rect 162814 667898 162986 668134
rect 163222 667898 163394 668134
rect 162814 632454 163394 667898
rect 162814 632218 162986 632454
rect 163222 632218 163394 632454
rect 162814 632134 163394 632218
rect 162814 631898 162986 632134
rect 163222 631898 163394 632134
rect 162814 596454 163394 631898
rect 162814 596218 162986 596454
rect 163222 596218 163394 596454
rect 162814 596134 163394 596218
rect 162814 595898 162986 596134
rect 163222 595898 163394 596134
rect 162814 560454 163394 595898
rect 162814 560218 162986 560454
rect 163222 560218 163394 560454
rect 162814 560134 163394 560218
rect 162814 559898 162986 560134
rect 163222 559898 163394 560134
rect 162814 524454 163394 559898
rect 162814 524218 162986 524454
rect 163222 524218 163394 524454
rect 162814 524134 163394 524218
rect 162814 523898 162986 524134
rect 163222 523898 163394 524134
rect 162814 488454 163394 523898
rect 162814 488218 162986 488454
rect 163222 488218 163394 488454
rect 162814 488134 163394 488218
rect 162814 487898 162986 488134
rect 163222 487898 163394 488134
rect 162814 452454 163394 487898
rect 162814 452218 162986 452454
rect 163222 452218 163394 452454
rect 162814 452134 163394 452218
rect 162814 451898 162986 452134
rect 163222 451898 163394 452134
rect 162814 416454 163394 451898
rect 162814 416218 162986 416454
rect 163222 416218 163394 416454
rect 162814 416134 163394 416218
rect 162814 415898 162986 416134
rect 163222 415898 163394 416134
rect 162814 380454 163394 415898
rect 162814 380218 162986 380454
rect 163222 380218 163394 380454
rect 162814 380134 163394 380218
rect 162814 379898 162986 380134
rect 163222 379898 163394 380134
rect 162814 344454 163394 379898
rect 162814 344218 162986 344454
rect 163222 344218 163394 344454
rect 162814 344134 163394 344218
rect 162814 343898 162986 344134
rect 163222 343898 163394 344134
rect 162814 308454 163394 343898
rect 162814 308218 162986 308454
rect 163222 308218 163394 308454
rect 162814 308134 163394 308218
rect 162814 307898 162986 308134
rect 163222 307898 163394 308134
rect 162814 272454 163394 307898
rect 162814 272218 162986 272454
rect 163222 272218 163394 272454
rect 162814 272134 163394 272218
rect 162814 271898 162986 272134
rect 163222 271898 163394 272134
rect 162814 236454 163394 271898
rect 162814 236218 162986 236454
rect 163222 236218 163394 236454
rect 162814 236134 163394 236218
rect 162814 235898 162986 236134
rect 163222 235898 163394 236134
rect 162814 200454 163394 235898
rect 162814 200218 162986 200454
rect 163222 200218 163394 200454
rect 162814 200134 163394 200218
rect 162814 199898 162986 200134
rect 163222 199898 163394 200134
rect 162814 164454 163394 199898
rect 162814 164218 162986 164454
rect 163222 164218 163394 164454
rect 162814 164134 163394 164218
rect 162814 163898 162986 164134
rect 163222 163898 163394 164134
rect 162814 128454 163394 163898
rect 162814 128218 162986 128454
rect 163222 128218 163394 128454
rect 162814 128134 163394 128218
rect 162814 127898 162986 128134
rect 163222 127898 163394 128134
rect 162814 92454 163394 127898
rect 162814 92218 162986 92454
rect 163222 92218 163394 92454
rect 162814 92134 163394 92218
rect 162814 91898 162986 92134
rect 163222 91898 163394 92134
rect 162814 56454 163394 91898
rect 162814 56218 162986 56454
rect 163222 56218 163394 56454
rect 162814 56134 163394 56218
rect 162814 55898 162986 56134
rect 163222 55898 163394 56134
rect 162814 20454 163394 55898
rect 162814 20218 162986 20454
rect 163222 20218 163394 20454
rect 162814 20134 163394 20218
rect 162814 19898 162986 20134
rect 163222 19898 163394 20134
rect 162814 -1266 163394 19898
rect 162814 -1502 162986 -1266
rect 163222 -1502 163394 -1266
rect 162814 -1586 163394 -1502
rect 162814 -1822 162986 -1586
rect 163222 -1822 163394 -1586
rect 162814 -1834 163394 -1822
rect 166294 671934 166874 707042
rect 166294 671698 166466 671934
rect 166702 671698 166874 671934
rect 166294 671614 166874 671698
rect 166294 671378 166466 671614
rect 166702 671378 166874 671614
rect 166294 635934 166874 671378
rect 166294 635698 166466 635934
rect 166702 635698 166874 635934
rect 166294 635614 166874 635698
rect 166294 635378 166466 635614
rect 166702 635378 166874 635614
rect 166294 599934 166874 635378
rect 166294 599698 166466 599934
rect 166702 599698 166874 599934
rect 166294 599614 166874 599698
rect 166294 599378 166466 599614
rect 166702 599378 166874 599614
rect 166294 563934 166874 599378
rect 166294 563698 166466 563934
rect 166702 563698 166874 563934
rect 166294 563614 166874 563698
rect 166294 563378 166466 563614
rect 166702 563378 166874 563614
rect 166294 527934 166874 563378
rect 166294 527698 166466 527934
rect 166702 527698 166874 527934
rect 166294 527614 166874 527698
rect 166294 527378 166466 527614
rect 166702 527378 166874 527614
rect 166294 491934 166874 527378
rect 166294 491698 166466 491934
rect 166702 491698 166874 491934
rect 166294 491614 166874 491698
rect 166294 491378 166466 491614
rect 166702 491378 166874 491614
rect 166294 455934 166874 491378
rect 166294 455698 166466 455934
rect 166702 455698 166874 455934
rect 166294 455614 166874 455698
rect 166294 455378 166466 455614
rect 166702 455378 166874 455614
rect 166294 419934 166874 455378
rect 166294 419698 166466 419934
rect 166702 419698 166874 419934
rect 166294 419614 166874 419698
rect 166294 419378 166466 419614
rect 166702 419378 166874 419614
rect 166294 383934 166874 419378
rect 166294 383698 166466 383934
rect 166702 383698 166874 383934
rect 166294 383614 166874 383698
rect 166294 383378 166466 383614
rect 166702 383378 166874 383614
rect 166294 347934 166874 383378
rect 166294 347698 166466 347934
rect 166702 347698 166874 347934
rect 166294 347614 166874 347698
rect 166294 347378 166466 347614
rect 166702 347378 166874 347614
rect 166294 311934 166874 347378
rect 166294 311698 166466 311934
rect 166702 311698 166874 311934
rect 166294 311614 166874 311698
rect 166294 311378 166466 311614
rect 166702 311378 166874 311614
rect 166294 275934 166874 311378
rect 166294 275698 166466 275934
rect 166702 275698 166874 275934
rect 166294 275614 166874 275698
rect 166294 275378 166466 275614
rect 166702 275378 166874 275614
rect 166294 239934 166874 275378
rect 166294 239698 166466 239934
rect 166702 239698 166874 239934
rect 166294 239614 166874 239698
rect 166294 239378 166466 239614
rect 166702 239378 166874 239614
rect 166294 203934 166874 239378
rect 166294 203698 166466 203934
rect 166702 203698 166874 203934
rect 166294 203614 166874 203698
rect 166294 203378 166466 203614
rect 166702 203378 166874 203614
rect 166294 167934 166874 203378
rect 166294 167698 166466 167934
rect 166702 167698 166874 167934
rect 166294 167614 166874 167698
rect 166294 167378 166466 167614
rect 166702 167378 166874 167614
rect 166294 131934 166874 167378
rect 166294 131698 166466 131934
rect 166702 131698 166874 131934
rect 166294 131614 166874 131698
rect 166294 131378 166466 131614
rect 166702 131378 166874 131614
rect 166294 95934 166874 131378
rect 166294 95698 166466 95934
rect 166702 95698 166874 95934
rect 166294 95614 166874 95698
rect 166294 95378 166466 95614
rect 166702 95378 166874 95614
rect 166294 59934 166874 95378
rect 166294 59698 166466 59934
rect 166702 59698 166874 59934
rect 166294 59614 166874 59698
rect 166294 59378 166466 59614
rect 166702 59378 166874 59614
rect 166294 23934 166874 59378
rect 166294 23698 166466 23934
rect 166702 23698 166874 23934
rect 166294 23614 166874 23698
rect 166294 23378 166466 23614
rect 166702 23378 166874 23614
rect 166294 -3106 166874 23378
rect 166294 -3342 166466 -3106
rect 166702 -3342 166874 -3106
rect 166294 -3426 166874 -3342
rect 166294 -3662 166466 -3426
rect 166702 -3662 166874 -3426
rect 166294 -3674 166874 -3662
rect 169774 675414 170354 708882
rect 169774 675178 169946 675414
rect 170182 675178 170354 675414
rect 169774 675094 170354 675178
rect 169774 674858 169946 675094
rect 170182 674858 170354 675094
rect 169774 639414 170354 674858
rect 169774 639178 169946 639414
rect 170182 639178 170354 639414
rect 169774 639094 170354 639178
rect 169774 638858 169946 639094
rect 170182 638858 170354 639094
rect 169774 603414 170354 638858
rect 169774 603178 169946 603414
rect 170182 603178 170354 603414
rect 169774 603094 170354 603178
rect 169774 602858 169946 603094
rect 170182 602858 170354 603094
rect 169774 567414 170354 602858
rect 169774 567178 169946 567414
rect 170182 567178 170354 567414
rect 169774 567094 170354 567178
rect 169774 566858 169946 567094
rect 170182 566858 170354 567094
rect 169774 531414 170354 566858
rect 169774 531178 169946 531414
rect 170182 531178 170354 531414
rect 169774 531094 170354 531178
rect 169774 530858 169946 531094
rect 170182 530858 170354 531094
rect 169774 495414 170354 530858
rect 169774 495178 169946 495414
rect 170182 495178 170354 495414
rect 169774 495094 170354 495178
rect 169774 494858 169946 495094
rect 170182 494858 170354 495094
rect 169774 459414 170354 494858
rect 169774 459178 169946 459414
rect 170182 459178 170354 459414
rect 169774 459094 170354 459178
rect 169774 458858 169946 459094
rect 170182 458858 170354 459094
rect 169774 423414 170354 458858
rect 169774 423178 169946 423414
rect 170182 423178 170354 423414
rect 169774 423094 170354 423178
rect 169774 422858 169946 423094
rect 170182 422858 170354 423094
rect 169774 387414 170354 422858
rect 169774 387178 169946 387414
rect 170182 387178 170354 387414
rect 169774 387094 170354 387178
rect 169774 386858 169946 387094
rect 170182 386858 170354 387094
rect 169774 351414 170354 386858
rect 169774 351178 169946 351414
rect 170182 351178 170354 351414
rect 169774 351094 170354 351178
rect 169774 350858 169946 351094
rect 170182 350858 170354 351094
rect 169774 315414 170354 350858
rect 169774 315178 169946 315414
rect 170182 315178 170354 315414
rect 169774 315094 170354 315178
rect 169774 314858 169946 315094
rect 170182 314858 170354 315094
rect 169774 279414 170354 314858
rect 169774 279178 169946 279414
rect 170182 279178 170354 279414
rect 169774 279094 170354 279178
rect 169774 278858 169946 279094
rect 170182 278858 170354 279094
rect 169774 243414 170354 278858
rect 169774 243178 169946 243414
rect 170182 243178 170354 243414
rect 169774 243094 170354 243178
rect 169774 242858 169946 243094
rect 170182 242858 170354 243094
rect 169774 207414 170354 242858
rect 169774 207178 169946 207414
rect 170182 207178 170354 207414
rect 169774 207094 170354 207178
rect 169774 206858 169946 207094
rect 170182 206858 170354 207094
rect 169774 171414 170354 206858
rect 169774 171178 169946 171414
rect 170182 171178 170354 171414
rect 169774 171094 170354 171178
rect 169774 170858 169946 171094
rect 170182 170858 170354 171094
rect 169774 135414 170354 170858
rect 169774 135178 169946 135414
rect 170182 135178 170354 135414
rect 169774 135094 170354 135178
rect 169774 134858 169946 135094
rect 170182 134858 170354 135094
rect 169774 99414 170354 134858
rect 169774 99178 169946 99414
rect 170182 99178 170354 99414
rect 169774 99094 170354 99178
rect 169774 98858 169946 99094
rect 170182 98858 170354 99094
rect 169774 63414 170354 98858
rect 169774 63178 169946 63414
rect 170182 63178 170354 63414
rect 169774 63094 170354 63178
rect 169774 62858 169946 63094
rect 170182 62858 170354 63094
rect 169774 27414 170354 62858
rect 169774 27178 169946 27414
rect 170182 27178 170354 27414
rect 169774 27094 170354 27178
rect 169774 26858 169946 27094
rect 170182 26858 170354 27094
rect 169774 -4946 170354 26858
rect 169774 -5182 169946 -4946
rect 170182 -5182 170354 -4946
rect 169774 -5266 170354 -5182
rect 169774 -5502 169946 -5266
rect 170182 -5502 170354 -5266
rect 169774 -5514 170354 -5502
rect 173254 678894 173834 710722
rect 191254 710358 191834 711290
rect 191254 710122 191426 710358
rect 191662 710122 191834 710358
rect 191254 710038 191834 710122
rect 191254 709802 191426 710038
rect 191662 709802 191834 710038
rect 187774 708518 188354 709450
rect 187774 708282 187946 708518
rect 188182 708282 188354 708518
rect 187774 708198 188354 708282
rect 187774 707962 187946 708198
rect 188182 707962 188354 708198
rect 184294 706678 184874 707610
rect 184294 706442 184466 706678
rect 184702 706442 184874 706678
rect 184294 706358 184874 706442
rect 184294 706122 184466 706358
rect 184702 706122 184874 706358
rect 173254 678658 173426 678894
rect 173662 678658 173834 678894
rect 173254 678574 173834 678658
rect 173254 678338 173426 678574
rect 173662 678338 173834 678574
rect 173254 642894 173834 678338
rect 173254 642658 173426 642894
rect 173662 642658 173834 642894
rect 173254 642574 173834 642658
rect 173254 642338 173426 642574
rect 173662 642338 173834 642574
rect 173254 606894 173834 642338
rect 173254 606658 173426 606894
rect 173662 606658 173834 606894
rect 173254 606574 173834 606658
rect 173254 606338 173426 606574
rect 173662 606338 173834 606574
rect 173254 570894 173834 606338
rect 173254 570658 173426 570894
rect 173662 570658 173834 570894
rect 173254 570574 173834 570658
rect 173254 570338 173426 570574
rect 173662 570338 173834 570574
rect 173254 534894 173834 570338
rect 173254 534658 173426 534894
rect 173662 534658 173834 534894
rect 173254 534574 173834 534658
rect 173254 534338 173426 534574
rect 173662 534338 173834 534574
rect 173254 498894 173834 534338
rect 173254 498658 173426 498894
rect 173662 498658 173834 498894
rect 173254 498574 173834 498658
rect 173254 498338 173426 498574
rect 173662 498338 173834 498574
rect 173254 462894 173834 498338
rect 173254 462658 173426 462894
rect 173662 462658 173834 462894
rect 173254 462574 173834 462658
rect 173254 462338 173426 462574
rect 173662 462338 173834 462574
rect 173254 426894 173834 462338
rect 173254 426658 173426 426894
rect 173662 426658 173834 426894
rect 173254 426574 173834 426658
rect 173254 426338 173426 426574
rect 173662 426338 173834 426574
rect 173254 390894 173834 426338
rect 173254 390658 173426 390894
rect 173662 390658 173834 390894
rect 173254 390574 173834 390658
rect 173254 390338 173426 390574
rect 173662 390338 173834 390574
rect 173254 354894 173834 390338
rect 173254 354658 173426 354894
rect 173662 354658 173834 354894
rect 173254 354574 173834 354658
rect 173254 354338 173426 354574
rect 173662 354338 173834 354574
rect 173254 318894 173834 354338
rect 173254 318658 173426 318894
rect 173662 318658 173834 318894
rect 173254 318574 173834 318658
rect 173254 318338 173426 318574
rect 173662 318338 173834 318574
rect 173254 282894 173834 318338
rect 173254 282658 173426 282894
rect 173662 282658 173834 282894
rect 173254 282574 173834 282658
rect 173254 282338 173426 282574
rect 173662 282338 173834 282574
rect 173254 246894 173834 282338
rect 173254 246658 173426 246894
rect 173662 246658 173834 246894
rect 173254 246574 173834 246658
rect 173254 246338 173426 246574
rect 173662 246338 173834 246574
rect 173254 210894 173834 246338
rect 173254 210658 173426 210894
rect 173662 210658 173834 210894
rect 173254 210574 173834 210658
rect 173254 210338 173426 210574
rect 173662 210338 173834 210574
rect 173254 174894 173834 210338
rect 173254 174658 173426 174894
rect 173662 174658 173834 174894
rect 173254 174574 173834 174658
rect 173254 174338 173426 174574
rect 173662 174338 173834 174574
rect 173254 138894 173834 174338
rect 173254 138658 173426 138894
rect 173662 138658 173834 138894
rect 173254 138574 173834 138658
rect 173254 138338 173426 138574
rect 173662 138338 173834 138574
rect 173254 102894 173834 138338
rect 173254 102658 173426 102894
rect 173662 102658 173834 102894
rect 173254 102574 173834 102658
rect 173254 102338 173426 102574
rect 173662 102338 173834 102574
rect 173254 66894 173834 102338
rect 173254 66658 173426 66894
rect 173662 66658 173834 66894
rect 173254 66574 173834 66658
rect 173254 66338 173426 66574
rect 173662 66338 173834 66574
rect 173254 30894 173834 66338
rect 173254 30658 173426 30894
rect 173662 30658 173834 30894
rect 173254 30574 173834 30658
rect 173254 30338 173426 30574
rect 173662 30338 173834 30574
rect 155254 -6102 155426 -5866
rect 155662 -6102 155834 -5866
rect 155254 -6186 155834 -6102
rect 155254 -6422 155426 -6186
rect 155662 -6422 155834 -6186
rect 155254 -7354 155834 -6422
rect 173254 -6786 173834 30338
rect 180814 704838 181394 705770
rect 180814 704602 180986 704838
rect 181222 704602 181394 704838
rect 180814 704518 181394 704602
rect 180814 704282 180986 704518
rect 181222 704282 181394 704518
rect 180814 686454 181394 704282
rect 180814 686218 180986 686454
rect 181222 686218 181394 686454
rect 180814 686134 181394 686218
rect 180814 685898 180986 686134
rect 181222 685898 181394 686134
rect 180814 650454 181394 685898
rect 180814 650218 180986 650454
rect 181222 650218 181394 650454
rect 180814 650134 181394 650218
rect 180814 649898 180986 650134
rect 181222 649898 181394 650134
rect 180814 614454 181394 649898
rect 180814 614218 180986 614454
rect 181222 614218 181394 614454
rect 180814 614134 181394 614218
rect 180814 613898 180986 614134
rect 181222 613898 181394 614134
rect 180814 578454 181394 613898
rect 180814 578218 180986 578454
rect 181222 578218 181394 578454
rect 180814 578134 181394 578218
rect 180814 577898 180986 578134
rect 181222 577898 181394 578134
rect 180814 542454 181394 577898
rect 180814 542218 180986 542454
rect 181222 542218 181394 542454
rect 180814 542134 181394 542218
rect 180814 541898 180986 542134
rect 181222 541898 181394 542134
rect 180814 506454 181394 541898
rect 180814 506218 180986 506454
rect 181222 506218 181394 506454
rect 180814 506134 181394 506218
rect 180814 505898 180986 506134
rect 181222 505898 181394 506134
rect 180814 470454 181394 505898
rect 180814 470218 180986 470454
rect 181222 470218 181394 470454
rect 180814 470134 181394 470218
rect 180814 469898 180986 470134
rect 181222 469898 181394 470134
rect 180814 434454 181394 469898
rect 180814 434218 180986 434454
rect 181222 434218 181394 434454
rect 180814 434134 181394 434218
rect 180814 433898 180986 434134
rect 181222 433898 181394 434134
rect 180814 398454 181394 433898
rect 180814 398218 180986 398454
rect 181222 398218 181394 398454
rect 180814 398134 181394 398218
rect 180814 397898 180986 398134
rect 181222 397898 181394 398134
rect 180814 362454 181394 397898
rect 180814 362218 180986 362454
rect 181222 362218 181394 362454
rect 180814 362134 181394 362218
rect 180814 361898 180986 362134
rect 181222 361898 181394 362134
rect 180814 326454 181394 361898
rect 180814 326218 180986 326454
rect 181222 326218 181394 326454
rect 180814 326134 181394 326218
rect 180814 325898 180986 326134
rect 181222 325898 181394 326134
rect 180814 290454 181394 325898
rect 180814 290218 180986 290454
rect 181222 290218 181394 290454
rect 180814 290134 181394 290218
rect 180814 289898 180986 290134
rect 181222 289898 181394 290134
rect 180814 254454 181394 289898
rect 180814 254218 180986 254454
rect 181222 254218 181394 254454
rect 180814 254134 181394 254218
rect 180814 253898 180986 254134
rect 181222 253898 181394 254134
rect 180814 218454 181394 253898
rect 180814 218218 180986 218454
rect 181222 218218 181394 218454
rect 180814 218134 181394 218218
rect 180814 217898 180986 218134
rect 181222 217898 181394 218134
rect 180814 182454 181394 217898
rect 180814 182218 180986 182454
rect 181222 182218 181394 182454
rect 180814 182134 181394 182218
rect 180814 181898 180986 182134
rect 181222 181898 181394 182134
rect 180814 146454 181394 181898
rect 180814 146218 180986 146454
rect 181222 146218 181394 146454
rect 180814 146134 181394 146218
rect 180814 145898 180986 146134
rect 181222 145898 181394 146134
rect 180814 110454 181394 145898
rect 180814 110218 180986 110454
rect 181222 110218 181394 110454
rect 180814 110134 181394 110218
rect 180814 109898 180986 110134
rect 181222 109898 181394 110134
rect 180814 74454 181394 109898
rect 180814 74218 180986 74454
rect 181222 74218 181394 74454
rect 180814 74134 181394 74218
rect 180814 73898 180986 74134
rect 181222 73898 181394 74134
rect 180814 38454 181394 73898
rect 180814 38218 180986 38454
rect 181222 38218 181394 38454
rect 180814 38134 181394 38218
rect 180814 37898 180986 38134
rect 181222 37898 181394 38134
rect 180814 2454 181394 37898
rect 180814 2218 180986 2454
rect 181222 2218 181394 2454
rect 180814 2134 181394 2218
rect 180814 1898 180986 2134
rect 181222 1898 181394 2134
rect 180814 -346 181394 1898
rect 180814 -582 180986 -346
rect 181222 -582 181394 -346
rect 180814 -666 181394 -582
rect 180814 -902 180986 -666
rect 181222 -902 181394 -666
rect 180814 -1834 181394 -902
rect 184294 689934 184874 706122
rect 184294 689698 184466 689934
rect 184702 689698 184874 689934
rect 184294 689614 184874 689698
rect 184294 689378 184466 689614
rect 184702 689378 184874 689614
rect 184294 653934 184874 689378
rect 184294 653698 184466 653934
rect 184702 653698 184874 653934
rect 184294 653614 184874 653698
rect 184294 653378 184466 653614
rect 184702 653378 184874 653614
rect 184294 617934 184874 653378
rect 184294 617698 184466 617934
rect 184702 617698 184874 617934
rect 184294 617614 184874 617698
rect 184294 617378 184466 617614
rect 184702 617378 184874 617614
rect 184294 581934 184874 617378
rect 184294 581698 184466 581934
rect 184702 581698 184874 581934
rect 184294 581614 184874 581698
rect 184294 581378 184466 581614
rect 184702 581378 184874 581614
rect 184294 545934 184874 581378
rect 184294 545698 184466 545934
rect 184702 545698 184874 545934
rect 184294 545614 184874 545698
rect 184294 545378 184466 545614
rect 184702 545378 184874 545614
rect 184294 509934 184874 545378
rect 184294 509698 184466 509934
rect 184702 509698 184874 509934
rect 184294 509614 184874 509698
rect 184294 509378 184466 509614
rect 184702 509378 184874 509614
rect 184294 473934 184874 509378
rect 184294 473698 184466 473934
rect 184702 473698 184874 473934
rect 184294 473614 184874 473698
rect 184294 473378 184466 473614
rect 184702 473378 184874 473614
rect 184294 437934 184874 473378
rect 184294 437698 184466 437934
rect 184702 437698 184874 437934
rect 184294 437614 184874 437698
rect 184294 437378 184466 437614
rect 184702 437378 184874 437614
rect 184294 401934 184874 437378
rect 184294 401698 184466 401934
rect 184702 401698 184874 401934
rect 184294 401614 184874 401698
rect 184294 401378 184466 401614
rect 184702 401378 184874 401614
rect 184294 365934 184874 401378
rect 184294 365698 184466 365934
rect 184702 365698 184874 365934
rect 184294 365614 184874 365698
rect 184294 365378 184466 365614
rect 184702 365378 184874 365614
rect 184294 329934 184874 365378
rect 184294 329698 184466 329934
rect 184702 329698 184874 329934
rect 184294 329614 184874 329698
rect 184294 329378 184466 329614
rect 184702 329378 184874 329614
rect 184294 293934 184874 329378
rect 184294 293698 184466 293934
rect 184702 293698 184874 293934
rect 184294 293614 184874 293698
rect 184294 293378 184466 293614
rect 184702 293378 184874 293614
rect 184294 257934 184874 293378
rect 184294 257698 184466 257934
rect 184702 257698 184874 257934
rect 184294 257614 184874 257698
rect 184294 257378 184466 257614
rect 184702 257378 184874 257614
rect 184294 221934 184874 257378
rect 184294 221698 184466 221934
rect 184702 221698 184874 221934
rect 184294 221614 184874 221698
rect 184294 221378 184466 221614
rect 184702 221378 184874 221614
rect 184294 185934 184874 221378
rect 184294 185698 184466 185934
rect 184702 185698 184874 185934
rect 184294 185614 184874 185698
rect 184294 185378 184466 185614
rect 184702 185378 184874 185614
rect 184294 149934 184874 185378
rect 184294 149698 184466 149934
rect 184702 149698 184874 149934
rect 184294 149614 184874 149698
rect 184294 149378 184466 149614
rect 184702 149378 184874 149614
rect 184294 113934 184874 149378
rect 184294 113698 184466 113934
rect 184702 113698 184874 113934
rect 184294 113614 184874 113698
rect 184294 113378 184466 113614
rect 184702 113378 184874 113614
rect 184294 77934 184874 113378
rect 184294 77698 184466 77934
rect 184702 77698 184874 77934
rect 184294 77614 184874 77698
rect 184294 77378 184466 77614
rect 184702 77378 184874 77614
rect 184294 41934 184874 77378
rect 184294 41698 184466 41934
rect 184702 41698 184874 41934
rect 184294 41614 184874 41698
rect 184294 41378 184466 41614
rect 184702 41378 184874 41614
rect 184294 5934 184874 41378
rect 184294 5698 184466 5934
rect 184702 5698 184874 5934
rect 184294 5614 184874 5698
rect 184294 5378 184466 5614
rect 184702 5378 184874 5614
rect 184294 -2186 184874 5378
rect 184294 -2422 184466 -2186
rect 184702 -2422 184874 -2186
rect 184294 -2506 184874 -2422
rect 184294 -2742 184466 -2506
rect 184702 -2742 184874 -2506
rect 184294 -3674 184874 -2742
rect 187774 693414 188354 707962
rect 187774 693178 187946 693414
rect 188182 693178 188354 693414
rect 187774 693094 188354 693178
rect 187774 692858 187946 693094
rect 188182 692858 188354 693094
rect 187774 657414 188354 692858
rect 187774 657178 187946 657414
rect 188182 657178 188354 657414
rect 187774 657094 188354 657178
rect 187774 656858 187946 657094
rect 188182 656858 188354 657094
rect 187774 621414 188354 656858
rect 187774 621178 187946 621414
rect 188182 621178 188354 621414
rect 187774 621094 188354 621178
rect 187774 620858 187946 621094
rect 188182 620858 188354 621094
rect 187774 585414 188354 620858
rect 187774 585178 187946 585414
rect 188182 585178 188354 585414
rect 187774 585094 188354 585178
rect 187774 584858 187946 585094
rect 188182 584858 188354 585094
rect 187774 549414 188354 584858
rect 187774 549178 187946 549414
rect 188182 549178 188354 549414
rect 187774 549094 188354 549178
rect 187774 548858 187946 549094
rect 188182 548858 188354 549094
rect 187774 513414 188354 548858
rect 187774 513178 187946 513414
rect 188182 513178 188354 513414
rect 187774 513094 188354 513178
rect 187774 512858 187946 513094
rect 188182 512858 188354 513094
rect 187774 477414 188354 512858
rect 187774 477178 187946 477414
rect 188182 477178 188354 477414
rect 187774 477094 188354 477178
rect 187774 476858 187946 477094
rect 188182 476858 188354 477094
rect 187774 441414 188354 476858
rect 187774 441178 187946 441414
rect 188182 441178 188354 441414
rect 187774 441094 188354 441178
rect 187774 440858 187946 441094
rect 188182 440858 188354 441094
rect 187774 405414 188354 440858
rect 187774 405178 187946 405414
rect 188182 405178 188354 405414
rect 187774 405094 188354 405178
rect 187774 404858 187946 405094
rect 188182 404858 188354 405094
rect 187774 369414 188354 404858
rect 187774 369178 187946 369414
rect 188182 369178 188354 369414
rect 187774 369094 188354 369178
rect 187774 368858 187946 369094
rect 188182 368858 188354 369094
rect 187774 333414 188354 368858
rect 187774 333178 187946 333414
rect 188182 333178 188354 333414
rect 187774 333094 188354 333178
rect 187774 332858 187946 333094
rect 188182 332858 188354 333094
rect 187774 297414 188354 332858
rect 187774 297178 187946 297414
rect 188182 297178 188354 297414
rect 187774 297094 188354 297178
rect 187774 296858 187946 297094
rect 188182 296858 188354 297094
rect 187774 261414 188354 296858
rect 187774 261178 187946 261414
rect 188182 261178 188354 261414
rect 187774 261094 188354 261178
rect 187774 260858 187946 261094
rect 188182 260858 188354 261094
rect 187774 225414 188354 260858
rect 187774 225178 187946 225414
rect 188182 225178 188354 225414
rect 187774 225094 188354 225178
rect 187774 224858 187946 225094
rect 188182 224858 188354 225094
rect 187774 189414 188354 224858
rect 187774 189178 187946 189414
rect 188182 189178 188354 189414
rect 187774 189094 188354 189178
rect 187774 188858 187946 189094
rect 188182 188858 188354 189094
rect 187774 153414 188354 188858
rect 187774 153178 187946 153414
rect 188182 153178 188354 153414
rect 187774 153094 188354 153178
rect 187774 152858 187946 153094
rect 188182 152858 188354 153094
rect 187774 117414 188354 152858
rect 187774 117178 187946 117414
rect 188182 117178 188354 117414
rect 187774 117094 188354 117178
rect 187774 116858 187946 117094
rect 188182 116858 188354 117094
rect 187774 81414 188354 116858
rect 187774 81178 187946 81414
rect 188182 81178 188354 81414
rect 187774 81094 188354 81178
rect 187774 80858 187946 81094
rect 188182 80858 188354 81094
rect 187774 45414 188354 80858
rect 187774 45178 187946 45414
rect 188182 45178 188354 45414
rect 187774 45094 188354 45178
rect 187774 44858 187946 45094
rect 188182 44858 188354 45094
rect 187774 9414 188354 44858
rect 187774 9178 187946 9414
rect 188182 9178 188354 9414
rect 187774 9094 188354 9178
rect 187774 8858 187946 9094
rect 188182 8858 188354 9094
rect 187774 -4026 188354 8858
rect 187774 -4262 187946 -4026
rect 188182 -4262 188354 -4026
rect 187774 -4346 188354 -4262
rect 187774 -4582 187946 -4346
rect 188182 -4582 188354 -4346
rect 187774 -5514 188354 -4582
rect 191254 696894 191834 709802
rect 209254 711278 209834 711290
rect 209254 711042 209426 711278
rect 209662 711042 209834 711278
rect 209254 710958 209834 711042
rect 209254 710722 209426 710958
rect 209662 710722 209834 710958
rect 205774 709438 206354 709450
rect 205774 709202 205946 709438
rect 206182 709202 206354 709438
rect 205774 709118 206354 709202
rect 205774 708882 205946 709118
rect 206182 708882 206354 709118
rect 202294 707598 202874 707610
rect 202294 707362 202466 707598
rect 202702 707362 202874 707598
rect 202294 707278 202874 707362
rect 202294 707042 202466 707278
rect 202702 707042 202874 707278
rect 191254 696658 191426 696894
rect 191662 696658 191834 696894
rect 191254 696574 191834 696658
rect 191254 696338 191426 696574
rect 191662 696338 191834 696574
rect 191254 660894 191834 696338
rect 191254 660658 191426 660894
rect 191662 660658 191834 660894
rect 191254 660574 191834 660658
rect 191254 660338 191426 660574
rect 191662 660338 191834 660574
rect 191254 624894 191834 660338
rect 191254 624658 191426 624894
rect 191662 624658 191834 624894
rect 191254 624574 191834 624658
rect 191254 624338 191426 624574
rect 191662 624338 191834 624574
rect 191254 588894 191834 624338
rect 191254 588658 191426 588894
rect 191662 588658 191834 588894
rect 191254 588574 191834 588658
rect 191254 588338 191426 588574
rect 191662 588338 191834 588574
rect 191254 552894 191834 588338
rect 191254 552658 191426 552894
rect 191662 552658 191834 552894
rect 191254 552574 191834 552658
rect 191254 552338 191426 552574
rect 191662 552338 191834 552574
rect 191254 516894 191834 552338
rect 191254 516658 191426 516894
rect 191662 516658 191834 516894
rect 191254 516574 191834 516658
rect 191254 516338 191426 516574
rect 191662 516338 191834 516574
rect 191254 480894 191834 516338
rect 191254 480658 191426 480894
rect 191662 480658 191834 480894
rect 191254 480574 191834 480658
rect 191254 480338 191426 480574
rect 191662 480338 191834 480574
rect 191254 444894 191834 480338
rect 191254 444658 191426 444894
rect 191662 444658 191834 444894
rect 191254 444574 191834 444658
rect 191254 444338 191426 444574
rect 191662 444338 191834 444574
rect 191254 408894 191834 444338
rect 191254 408658 191426 408894
rect 191662 408658 191834 408894
rect 191254 408574 191834 408658
rect 191254 408338 191426 408574
rect 191662 408338 191834 408574
rect 191254 372894 191834 408338
rect 191254 372658 191426 372894
rect 191662 372658 191834 372894
rect 191254 372574 191834 372658
rect 191254 372338 191426 372574
rect 191662 372338 191834 372574
rect 191254 336894 191834 372338
rect 191254 336658 191426 336894
rect 191662 336658 191834 336894
rect 191254 336574 191834 336658
rect 191254 336338 191426 336574
rect 191662 336338 191834 336574
rect 191254 300894 191834 336338
rect 191254 300658 191426 300894
rect 191662 300658 191834 300894
rect 191254 300574 191834 300658
rect 191254 300338 191426 300574
rect 191662 300338 191834 300574
rect 191254 264894 191834 300338
rect 191254 264658 191426 264894
rect 191662 264658 191834 264894
rect 191254 264574 191834 264658
rect 191254 264338 191426 264574
rect 191662 264338 191834 264574
rect 191254 228894 191834 264338
rect 191254 228658 191426 228894
rect 191662 228658 191834 228894
rect 191254 228574 191834 228658
rect 191254 228338 191426 228574
rect 191662 228338 191834 228574
rect 191254 192894 191834 228338
rect 191254 192658 191426 192894
rect 191662 192658 191834 192894
rect 191254 192574 191834 192658
rect 191254 192338 191426 192574
rect 191662 192338 191834 192574
rect 191254 156894 191834 192338
rect 191254 156658 191426 156894
rect 191662 156658 191834 156894
rect 191254 156574 191834 156658
rect 191254 156338 191426 156574
rect 191662 156338 191834 156574
rect 191254 120894 191834 156338
rect 191254 120658 191426 120894
rect 191662 120658 191834 120894
rect 191254 120574 191834 120658
rect 191254 120338 191426 120574
rect 191662 120338 191834 120574
rect 191254 84894 191834 120338
rect 191254 84658 191426 84894
rect 191662 84658 191834 84894
rect 191254 84574 191834 84658
rect 191254 84338 191426 84574
rect 191662 84338 191834 84574
rect 191254 48894 191834 84338
rect 191254 48658 191426 48894
rect 191662 48658 191834 48894
rect 191254 48574 191834 48658
rect 191254 48338 191426 48574
rect 191662 48338 191834 48574
rect 191254 12894 191834 48338
rect 191254 12658 191426 12894
rect 191662 12658 191834 12894
rect 191254 12574 191834 12658
rect 191254 12338 191426 12574
rect 191662 12338 191834 12574
rect 173254 -7022 173426 -6786
rect 173662 -7022 173834 -6786
rect 173254 -7106 173834 -7022
rect 173254 -7342 173426 -7106
rect 173662 -7342 173834 -7106
rect 173254 -7354 173834 -7342
rect 191254 -5866 191834 12338
rect 198814 705758 199394 705770
rect 198814 705522 198986 705758
rect 199222 705522 199394 705758
rect 198814 705438 199394 705522
rect 198814 705202 198986 705438
rect 199222 705202 199394 705438
rect 198814 668454 199394 705202
rect 198814 668218 198986 668454
rect 199222 668218 199394 668454
rect 198814 668134 199394 668218
rect 198814 667898 198986 668134
rect 199222 667898 199394 668134
rect 198814 632454 199394 667898
rect 198814 632218 198986 632454
rect 199222 632218 199394 632454
rect 198814 632134 199394 632218
rect 198814 631898 198986 632134
rect 199222 631898 199394 632134
rect 198814 596454 199394 631898
rect 198814 596218 198986 596454
rect 199222 596218 199394 596454
rect 198814 596134 199394 596218
rect 198814 595898 198986 596134
rect 199222 595898 199394 596134
rect 198814 560454 199394 595898
rect 198814 560218 198986 560454
rect 199222 560218 199394 560454
rect 198814 560134 199394 560218
rect 198814 559898 198986 560134
rect 199222 559898 199394 560134
rect 198814 524454 199394 559898
rect 198814 524218 198986 524454
rect 199222 524218 199394 524454
rect 198814 524134 199394 524218
rect 198814 523898 198986 524134
rect 199222 523898 199394 524134
rect 198814 488454 199394 523898
rect 198814 488218 198986 488454
rect 199222 488218 199394 488454
rect 198814 488134 199394 488218
rect 198814 487898 198986 488134
rect 199222 487898 199394 488134
rect 198814 452454 199394 487898
rect 198814 452218 198986 452454
rect 199222 452218 199394 452454
rect 198814 452134 199394 452218
rect 198814 451898 198986 452134
rect 199222 451898 199394 452134
rect 198814 416454 199394 451898
rect 198814 416218 198986 416454
rect 199222 416218 199394 416454
rect 198814 416134 199394 416218
rect 198814 415898 198986 416134
rect 199222 415898 199394 416134
rect 198814 380454 199394 415898
rect 198814 380218 198986 380454
rect 199222 380218 199394 380454
rect 198814 380134 199394 380218
rect 198814 379898 198986 380134
rect 199222 379898 199394 380134
rect 198814 344454 199394 379898
rect 198814 344218 198986 344454
rect 199222 344218 199394 344454
rect 198814 344134 199394 344218
rect 198814 343898 198986 344134
rect 199222 343898 199394 344134
rect 198814 308454 199394 343898
rect 198814 308218 198986 308454
rect 199222 308218 199394 308454
rect 198814 308134 199394 308218
rect 198814 307898 198986 308134
rect 199222 307898 199394 308134
rect 198814 272454 199394 307898
rect 198814 272218 198986 272454
rect 199222 272218 199394 272454
rect 198814 272134 199394 272218
rect 198814 271898 198986 272134
rect 199222 271898 199394 272134
rect 198814 236454 199394 271898
rect 198814 236218 198986 236454
rect 199222 236218 199394 236454
rect 198814 236134 199394 236218
rect 198814 235898 198986 236134
rect 199222 235898 199394 236134
rect 198814 200454 199394 235898
rect 198814 200218 198986 200454
rect 199222 200218 199394 200454
rect 198814 200134 199394 200218
rect 198814 199898 198986 200134
rect 199222 199898 199394 200134
rect 198814 164454 199394 199898
rect 198814 164218 198986 164454
rect 199222 164218 199394 164454
rect 198814 164134 199394 164218
rect 198814 163898 198986 164134
rect 199222 163898 199394 164134
rect 198814 128454 199394 163898
rect 198814 128218 198986 128454
rect 199222 128218 199394 128454
rect 198814 128134 199394 128218
rect 198814 127898 198986 128134
rect 199222 127898 199394 128134
rect 198814 92454 199394 127898
rect 198814 92218 198986 92454
rect 199222 92218 199394 92454
rect 198814 92134 199394 92218
rect 198814 91898 198986 92134
rect 199222 91898 199394 92134
rect 198814 56454 199394 91898
rect 198814 56218 198986 56454
rect 199222 56218 199394 56454
rect 198814 56134 199394 56218
rect 198814 55898 198986 56134
rect 199222 55898 199394 56134
rect 198814 20454 199394 55898
rect 198814 20218 198986 20454
rect 199222 20218 199394 20454
rect 198814 20134 199394 20218
rect 198814 19898 198986 20134
rect 199222 19898 199394 20134
rect 198814 -1266 199394 19898
rect 198814 -1502 198986 -1266
rect 199222 -1502 199394 -1266
rect 198814 -1586 199394 -1502
rect 198814 -1822 198986 -1586
rect 199222 -1822 199394 -1586
rect 198814 -1834 199394 -1822
rect 202294 671934 202874 707042
rect 202294 671698 202466 671934
rect 202702 671698 202874 671934
rect 202294 671614 202874 671698
rect 202294 671378 202466 671614
rect 202702 671378 202874 671614
rect 202294 635934 202874 671378
rect 202294 635698 202466 635934
rect 202702 635698 202874 635934
rect 202294 635614 202874 635698
rect 202294 635378 202466 635614
rect 202702 635378 202874 635614
rect 202294 599934 202874 635378
rect 202294 599698 202466 599934
rect 202702 599698 202874 599934
rect 202294 599614 202874 599698
rect 202294 599378 202466 599614
rect 202702 599378 202874 599614
rect 202294 563934 202874 599378
rect 202294 563698 202466 563934
rect 202702 563698 202874 563934
rect 202294 563614 202874 563698
rect 202294 563378 202466 563614
rect 202702 563378 202874 563614
rect 202294 527934 202874 563378
rect 202294 527698 202466 527934
rect 202702 527698 202874 527934
rect 202294 527614 202874 527698
rect 202294 527378 202466 527614
rect 202702 527378 202874 527614
rect 202294 491934 202874 527378
rect 202294 491698 202466 491934
rect 202702 491698 202874 491934
rect 202294 491614 202874 491698
rect 202294 491378 202466 491614
rect 202702 491378 202874 491614
rect 202294 455934 202874 491378
rect 202294 455698 202466 455934
rect 202702 455698 202874 455934
rect 202294 455614 202874 455698
rect 202294 455378 202466 455614
rect 202702 455378 202874 455614
rect 202294 419934 202874 455378
rect 202294 419698 202466 419934
rect 202702 419698 202874 419934
rect 202294 419614 202874 419698
rect 202294 419378 202466 419614
rect 202702 419378 202874 419614
rect 202294 383934 202874 419378
rect 202294 383698 202466 383934
rect 202702 383698 202874 383934
rect 202294 383614 202874 383698
rect 202294 383378 202466 383614
rect 202702 383378 202874 383614
rect 202294 347934 202874 383378
rect 202294 347698 202466 347934
rect 202702 347698 202874 347934
rect 202294 347614 202874 347698
rect 202294 347378 202466 347614
rect 202702 347378 202874 347614
rect 202294 311934 202874 347378
rect 202294 311698 202466 311934
rect 202702 311698 202874 311934
rect 202294 311614 202874 311698
rect 202294 311378 202466 311614
rect 202702 311378 202874 311614
rect 202294 275934 202874 311378
rect 202294 275698 202466 275934
rect 202702 275698 202874 275934
rect 202294 275614 202874 275698
rect 202294 275378 202466 275614
rect 202702 275378 202874 275614
rect 202294 239934 202874 275378
rect 202294 239698 202466 239934
rect 202702 239698 202874 239934
rect 202294 239614 202874 239698
rect 202294 239378 202466 239614
rect 202702 239378 202874 239614
rect 202294 203934 202874 239378
rect 202294 203698 202466 203934
rect 202702 203698 202874 203934
rect 202294 203614 202874 203698
rect 202294 203378 202466 203614
rect 202702 203378 202874 203614
rect 202294 167934 202874 203378
rect 202294 167698 202466 167934
rect 202702 167698 202874 167934
rect 202294 167614 202874 167698
rect 202294 167378 202466 167614
rect 202702 167378 202874 167614
rect 202294 131934 202874 167378
rect 202294 131698 202466 131934
rect 202702 131698 202874 131934
rect 202294 131614 202874 131698
rect 202294 131378 202466 131614
rect 202702 131378 202874 131614
rect 202294 95934 202874 131378
rect 202294 95698 202466 95934
rect 202702 95698 202874 95934
rect 202294 95614 202874 95698
rect 202294 95378 202466 95614
rect 202702 95378 202874 95614
rect 202294 59934 202874 95378
rect 202294 59698 202466 59934
rect 202702 59698 202874 59934
rect 202294 59614 202874 59698
rect 202294 59378 202466 59614
rect 202702 59378 202874 59614
rect 202294 23934 202874 59378
rect 202294 23698 202466 23934
rect 202702 23698 202874 23934
rect 202294 23614 202874 23698
rect 202294 23378 202466 23614
rect 202702 23378 202874 23614
rect 202294 -3106 202874 23378
rect 202294 -3342 202466 -3106
rect 202702 -3342 202874 -3106
rect 202294 -3426 202874 -3342
rect 202294 -3662 202466 -3426
rect 202702 -3662 202874 -3426
rect 202294 -3674 202874 -3662
rect 205774 675414 206354 708882
rect 205774 675178 205946 675414
rect 206182 675178 206354 675414
rect 205774 675094 206354 675178
rect 205774 674858 205946 675094
rect 206182 674858 206354 675094
rect 205774 639414 206354 674858
rect 205774 639178 205946 639414
rect 206182 639178 206354 639414
rect 205774 639094 206354 639178
rect 205774 638858 205946 639094
rect 206182 638858 206354 639094
rect 205774 603414 206354 638858
rect 205774 603178 205946 603414
rect 206182 603178 206354 603414
rect 205774 603094 206354 603178
rect 205774 602858 205946 603094
rect 206182 602858 206354 603094
rect 205774 567414 206354 602858
rect 205774 567178 205946 567414
rect 206182 567178 206354 567414
rect 205774 567094 206354 567178
rect 205774 566858 205946 567094
rect 206182 566858 206354 567094
rect 205774 531414 206354 566858
rect 205774 531178 205946 531414
rect 206182 531178 206354 531414
rect 205774 531094 206354 531178
rect 205774 530858 205946 531094
rect 206182 530858 206354 531094
rect 205774 495414 206354 530858
rect 205774 495178 205946 495414
rect 206182 495178 206354 495414
rect 205774 495094 206354 495178
rect 205774 494858 205946 495094
rect 206182 494858 206354 495094
rect 205774 459414 206354 494858
rect 205774 459178 205946 459414
rect 206182 459178 206354 459414
rect 205774 459094 206354 459178
rect 205774 458858 205946 459094
rect 206182 458858 206354 459094
rect 205774 423414 206354 458858
rect 205774 423178 205946 423414
rect 206182 423178 206354 423414
rect 205774 423094 206354 423178
rect 205774 422858 205946 423094
rect 206182 422858 206354 423094
rect 205774 387414 206354 422858
rect 205774 387178 205946 387414
rect 206182 387178 206354 387414
rect 205774 387094 206354 387178
rect 205774 386858 205946 387094
rect 206182 386858 206354 387094
rect 205774 351414 206354 386858
rect 205774 351178 205946 351414
rect 206182 351178 206354 351414
rect 205774 351094 206354 351178
rect 205774 350858 205946 351094
rect 206182 350858 206354 351094
rect 205774 315414 206354 350858
rect 205774 315178 205946 315414
rect 206182 315178 206354 315414
rect 205774 315094 206354 315178
rect 205774 314858 205946 315094
rect 206182 314858 206354 315094
rect 205774 279414 206354 314858
rect 205774 279178 205946 279414
rect 206182 279178 206354 279414
rect 205774 279094 206354 279178
rect 205774 278858 205946 279094
rect 206182 278858 206354 279094
rect 205774 243414 206354 278858
rect 205774 243178 205946 243414
rect 206182 243178 206354 243414
rect 205774 243094 206354 243178
rect 205774 242858 205946 243094
rect 206182 242858 206354 243094
rect 205774 207414 206354 242858
rect 205774 207178 205946 207414
rect 206182 207178 206354 207414
rect 205774 207094 206354 207178
rect 205774 206858 205946 207094
rect 206182 206858 206354 207094
rect 205774 171414 206354 206858
rect 205774 171178 205946 171414
rect 206182 171178 206354 171414
rect 205774 171094 206354 171178
rect 205774 170858 205946 171094
rect 206182 170858 206354 171094
rect 205774 135414 206354 170858
rect 205774 135178 205946 135414
rect 206182 135178 206354 135414
rect 205774 135094 206354 135178
rect 205774 134858 205946 135094
rect 206182 134858 206354 135094
rect 205774 99414 206354 134858
rect 205774 99178 205946 99414
rect 206182 99178 206354 99414
rect 205774 99094 206354 99178
rect 205774 98858 205946 99094
rect 206182 98858 206354 99094
rect 205774 63414 206354 98858
rect 205774 63178 205946 63414
rect 206182 63178 206354 63414
rect 205774 63094 206354 63178
rect 205774 62858 205946 63094
rect 206182 62858 206354 63094
rect 205774 27414 206354 62858
rect 205774 27178 205946 27414
rect 206182 27178 206354 27414
rect 205774 27094 206354 27178
rect 205774 26858 205946 27094
rect 206182 26858 206354 27094
rect 205774 -4946 206354 26858
rect 205774 -5182 205946 -4946
rect 206182 -5182 206354 -4946
rect 205774 -5266 206354 -5182
rect 205774 -5502 205946 -5266
rect 206182 -5502 206354 -5266
rect 205774 -5514 206354 -5502
rect 209254 678894 209834 710722
rect 227254 710358 227834 711290
rect 227254 710122 227426 710358
rect 227662 710122 227834 710358
rect 227254 710038 227834 710122
rect 227254 709802 227426 710038
rect 227662 709802 227834 710038
rect 223774 708518 224354 709450
rect 223774 708282 223946 708518
rect 224182 708282 224354 708518
rect 223774 708198 224354 708282
rect 223774 707962 223946 708198
rect 224182 707962 224354 708198
rect 220294 706678 220874 707610
rect 220294 706442 220466 706678
rect 220702 706442 220874 706678
rect 220294 706358 220874 706442
rect 220294 706122 220466 706358
rect 220702 706122 220874 706358
rect 209254 678658 209426 678894
rect 209662 678658 209834 678894
rect 209254 678574 209834 678658
rect 209254 678338 209426 678574
rect 209662 678338 209834 678574
rect 209254 642894 209834 678338
rect 209254 642658 209426 642894
rect 209662 642658 209834 642894
rect 209254 642574 209834 642658
rect 209254 642338 209426 642574
rect 209662 642338 209834 642574
rect 209254 606894 209834 642338
rect 209254 606658 209426 606894
rect 209662 606658 209834 606894
rect 209254 606574 209834 606658
rect 209254 606338 209426 606574
rect 209662 606338 209834 606574
rect 209254 570894 209834 606338
rect 209254 570658 209426 570894
rect 209662 570658 209834 570894
rect 209254 570574 209834 570658
rect 209254 570338 209426 570574
rect 209662 570338 209834 570574
rect 209254 534894 209834 570338
rect 209254 534658 209426 534894
rect 209662 534658 209834 534894
rect 209254 534574 209834 534658
rect 209254 534338 209426 534574
rect 209662 534338 209834 534574
rect 209254 498894 209834 534338
rect 209254 498658 209426 498894
rect 209662 498658 209834 498894
rect 209254 498574 209834 498658
rect 209254 498338 209426 498574
rect 209662 498338 209834 498574
rect 209254 462894 209834 498338
rect 209254 462658 209426 462894
rect 209662 462658 209834 462894
rect 209254 462574 209834 462658
rect 209254 462338 209426 462574
rect 209662 462338 209834 462574
rect 209254 426894 209834 462338
rect 209254 426658 209426 426894
rect 209662 426658 209834 426894
rect 209254 426574 209834 426658
rect 209254 426338 209426 426574
rect 209662 426338 209834 426574
rect 209254 390894 209834 426338
rect 209254 390658 209426 390894
rect 209662 390658 209834 390894
rect 209254 390574 209834 390658
rect 209254 390338 209426 390574
rect 209662 390338 209834 390574
rect 209254 354894 209834 390338
rect 209254 354658 209426 354894
rect 209662 354658 209834 354894
rect 209254 354574 209834 354658
rect 209254 354338 209426 354574
rect 209662 354338 209834 354574
rect 209254 318894 209834 354338
rect 209254 318658 209426 318894
rect 209662 318658 209834 318894
rect 209254 318574 209834 318658
rect 209254 318338 209426 318574
rect 209662 318338 209834 318574
rect 209254 282894 209834 318338
rect 209254 282658 209426 282894
rect 209662 282658 209834 282894
rect 209254 282574 209834 282658
rect 209254 282338 209426 282574
rect 209662 282338 209834 282574
rect 209254 246894 209834 282338
rect 209254 246658 209426 246894
rect 209662 246658 209834 246894
rect 209254 246574 209834 246658
rect 209254 246338 209426 246574
rect 209662 246338 209834 246574
rect 209254 210894 209834 246338
rect 209254 210658 209426 210894
rect 209662 210658 209834 210894
rect 209254 210574 209834 210658
rect 209254 210338 209426 210574
rect 209662 210338 209834 210574
rect 209254 174894 209834 210338
rect 209254 174658 209426 174894
rect 209662 174658 209834 174894
rect 209254 174574 209834 174658
rect 209254 174338 209426 174574
rect 209662 174338 209834 174574
rect 209254 138894 209834 174338
rect 209254 138658 209426 138894
rect 209662 138658 209834 138894
rect 209254 138574 209834 138658
rect 209254 138338 209426 138574
rect 209662 138338 209834 138574
rect 209254 102894 209834 138338
rect 209254 102658 209426 102894
rect 209662 102658 209834 102894
rect 209254 102574 209834 102658
rect 209254 102338 209426 102574
rect 209662 102338 209834 102574
rect 209254 66894 209834 102338
rect 209254 66658 209426 66894
rect 209662 66658 209834 66894
rect 209254 66574 209834 66658
rect 209254 66338 209426 66574
rect 209662 66338 209834 66574
rect 209254 30894 209834 66338
rect 209254 30658 209426 30894
rect 209662 30658 209834 30894
rect 209254 30574 209834 30658
rect 209254 30338 209426 30574
rect 209662 30338 209834 30574
rect 191254 -6102 191426 -5866
rect 191662 -6102 191834 -5866
rect 191254 -6186 191834 -6102
rect 191254 -6422 191426 -6186
rect 191662 -6422 191834 -6186
rect 191254 -7354 191834 -6422
rect 209254 -6786 209834 30338
rect 216814 704838 217394 705770
rect 216814 704602 216986 704838
rect 217222 704602 217394 704838
rect 216814 704518 217394 704602
rect 216814 704282 216986 704518
rect 217222 704282 217394 704518
rect 216814 686454 217394 704282
rect 216814 686218 216986 686454
rect 217222 686218 217394 686454
rect 216814 686134 217394 686218
rect 216814 685898 216986 686134
rect 217222 685898 217394 686134
rect 216814 650454 217394 685898
rect 216814 650218 216986 650454
rect 217222 650218 217394 650454
rect 216814 650134 217394 650218
rect 216814 649898 216986 650134
rect 217222 649898 217394 650134
rect 216814 614454 217394 649898
rect 216814 614218 216986 614454
rect 217222 614218 217394 614454
rect 216814 614134 217394 614218
rect 216814 613898 216986 614134
rect 217222 613898 217394 614134
rect 216814 578454 217394 613898
rect 216814 578218 216986 578454
rect 217222 578218 217394 578454
rect 216814 578134 217394 578218
rect 216814 577898 216986 578134
rect 217222 577898 217394 578134
rect 216814 542454 217394 577898
rect 216814 542218 216986 542454
rect 217222 542218 217394 542454
rect 216814 542134 217394 542218
rect 216814 541898 216986 542134
rect 217222 541898 217394 542134
rect 216814 506454 217394 541898
rect 216814 506218 216986 506454
rect 217222 506218 217394 506454
rect 216814 506134 217394 506218
rect 216814 505898 216986 506134
rect 217222 505898 217394 506134
rect 216814 470454 217394 505898
rect 216814 470218 216986 470454
rect 217222 470218 217394 470454
rect 216814 470134 217394 470218
rect 216814 469898 216986 470134
rect 217222 469898 217394 470134
rect 216814 434454 217394 469898
rect 216814 434218 216986 434454
rect 217222 434218 217394 434454
rect 216814 434134 217394 434218
rect 216814 433898 216986 434134
rect 217222 433898 217394 434134
rect 216814 398454 217394 433898
rect 216814 398218 216986 398454
rect 217222 398218 217394 398454
rect 216814 398134 217394 398218
rect 216814 397898 216986 398134
rect 217222 397898 217394 398134
rect 216814 362454 217394 397898
rect 216814 362218 216986 362454
rect 217222 362218 217394 362454
rect 216814 362134 217394 362218
rect 216814 361898 216986 362134
rect 217222 361898 217394 362134
rect 216814 326454 217394 361898
rect 216814 326218 216986 326454
rect 217222 326218 217394 326454
rect 216814 326134 217394 326218
rect 216814 325898 216986 326134
rect 217222 325898 217394 326134
rect 216814 290454 217394 325898
rect 216814 290218 216986 290454
rect 217222 290218 217394 290454
rect 216814 290134 217394 290218
rect 216814 289898 216986 290134
rect 217222 289898 217394 290134
rect 216814 254454 217394 289898
rect 216814 254218 216986 254454
rect 217222 254218 217394 254454
rect 216814 254134 217394 254218
rect 216814 253898 216986 254134
rect 217222 253898 217394 254134
rect 216814 218454 217394 253898
rect 216814 218218 216986 218454
rect 217222 218218 217394 218454
rect 216814 218134 217394 218218
rect 216814 217898 216986 218134
rect 217222 217898 217394 218134
rect 216814 182454 217394 217898
rect 216814 182218 216986 182454
rect 217222 182218 217394 182454
rect 216814 182134 217394 182218
rect 216814 181898 216986 182134
rect 217222 181898 217394 182134
rect 216814 146454 217394 181898
rect 216814 146218 216986 146454
rect 217222 146218 217394 146454
rect 216814 146134 217394 146218
rect 216814 145898 216986 146134
rect 217222 145898 217394 146134
rect 216814 110454 217394 145898
rect 216814 110218 216986 110454
rect 217222 110218 217394 110454
rect 216814 110134 217394 110218
rect 216814 109898 216986 110134
rect 217222 109898 217394 110134
rect 216814 74454 217394 109898
rect 216814 74218 216986 74454
rect 217222 74218 217394 74454
rect 216814 74134 217394 74218
rect 216814 73898 216986 74134
rect 217222 73898 217394 74134
rect 216814 38454 217394 73898
rect 216814 38218 216986 38454
rect 217222 38218 217394 38454
rect 216814 38134 217394 38218
rect 216814 37898 216986 38134
rect 217222 37898 217394 38134
rect 216814 2454 217394 37898
rect 216814 2218 216986 2454
rect 217222 2218 217394 2454
rect 216814 2134 217394 2218
rect 216814 1898 216986 2134
rect 217222 1898 217394 2134
rect 216814 -346 217394 1898
rect 216814 -582 216986 -346
rect 217222 -582 217394 -346
rect 216814 -666 217394 -582
rect 216814 -902 216986 -666
rect 217222 -902 217394 -666
rect 216814 -1834 217394 -902
rect 220294 689934 220874 706122
rect 220294 689698 220466 689934
rect 220702 689698 220874 689934
rect 220294 689614 220874 689698
rect 220294 689378 220466 689614
rect 220702 689378 220874 689614
rect 220294 653934 220874 689378
rect 220294 653698 220466 653934
rect 220702 653698 220874 653934
rect 220294 653614 220874 653698
rect 220294 653378 220466 653614
rect 220702 653378 220874 653614
rect 220294 617934 220874 653378
rect 220294 617698 220466 617934
rect 220702 617698 220874 617934
rect 220294 617614 220874 617698
rect 220294 617378 220466 617614
rect 220702 617378 220874 617614
rect 220294 581934 220874 617378
rect 220294 581698 220466 581934
rect 220702 581698 220874 581934
rect 220294 581614 220874 581698
rect 220294 581378 220466 581614
rect 220702 581378 220874 581614
rect 220294 545934 220874 581378
rect 220294 545698 220466 545934
rect 220702 545698 220874 545934
rect 220294 545614 220874 545698
rect 220294 545378 220466 545614
rect 220702 545378 220874 545614
rect 220294 509934 220874 545378
rect 220294 509698 220466 509934
rect 220702 509698 220874 509934
rect 220294 509614 220874 509698
rect 220294 509378 220466 509614
rect 220702 509378 220874 509614
rect 220294 473934 220874 509378
rect 220294 473698 220466 473934
rect 220702 473698 220874 473934
rect 220294 473614 220874 473698
rect 220294 473378 220466 473614
rect 220702 473378 220874 473614
rect 220294 437934 220874 473378
rect 220294 437698 220466 437934
rect 220702 437698 220874 437934
rect 220294 437614 220874 437698
rect 220294 437378 220466 437614
rect 220702 437378 220874 437614
rect 220294 401934 220874 437378
rect 220294 401698 220466 401934
rect 220702 401698 220874 401934
rect 220294 401614 220874 401698
rect 220294 401378 220466 401614
rect 220702 401378 220874 401614
rect 220294 365934 220874 401378
rect 220294 365698 220466 365934
rect 220702 365698 220874 365934
rect 220294 365614 220874 365698
rect 220294 365378 220466 365614
rect 220702 365378 220874 365614
rect 220294 329934 220874 365378
rect 220294 329698 220466 329934
rect 220702 329698 220874 329934
rect 220294 329614 220874 329698
rect 220294 329378 220466 329614
rect 220702 329378 220874 329614
rect 220294 293934 220874 329378
rect 220294 293698 220466 293934
rect 220702 293698 220874 293934
rect 220294 293614 220874 293698
rect 220294 293378 220466 293614
rect 220702 293378 220874 293614
rect 220294 257934 220874 293378
rect 220294 257698 220466 257934
rect 220702 257698 220874 257934
rect 220294 257614 220874 257698
rect 220294 257378 220466 257614
rect 220702 257378 220874 257614
rect 220294 221934 220874 257378
rect 220294 221698 220466 221934
rect 220702 221698 220874 221934
rect 220294 221614 220874 221698
rect 220294 221378 220466 221614
rect 220702 221378 220874 221614
rect 220294 185934 220874 221378
rect 220294 185698 220466 185934
rect 220702 185698 220874 185934
rect 220294 185614 220874 185698
rect 220294 185378 220466 185614
rect 220702 185378 220874 185614
rect 220294 149934 220874 185378
rect 220294 149698 220466 149934
rect 220702 149698 220874 149934
rect 220294 149614 220874 149698
rect 220294 149378 220466 149614
rect 220702 149378 220874 149614
rect 220294 113934 220874 149378
rect 220294 113698 220466 113934
rect 220702 113698 220874 113934
rect 220294 113614 220874 113698
rect 220294 113378 220466 113614
rect 220702 113378 220874 113614
rect 220294 77934 220874 113378
rect 220294 77698 220466 77934
rect 220702 77698 220874 77934
rect 220294 77614 220874 77698
rect 220294 77378 220466 77614
rect 220702 77378 220874 77614
rect 220294 41934 220874 77378
rect 220294 41698 220466 41934
rect 220702 41698 220874 41934
rect 220294 41614 220874 41698
rect 220294 41378 220466 41614
rect 220702 41378 220874 41614
rect 220294 5934 220874 41378
rect 220294 5698 220466 5934
rect 220702 5698 220874 5934
rect 220294 5614 220874 5698
rect 220294 5378 220466 5614
rect 220702 5378 220874 5614
rect 220294 -2186 220874 5378
rect 220294 -2422 220466 -2186
rect 220702 -2422 220874 -2186
rect 220294 -2506 220874 -2422
rect 220294 -2742 220466 -2506
rect 220702 -2742 220874 -2506
rect 220294 -3674 220874 -2742
rect 223774 693414 224354 707962
rect 223774 693178 223946 693414
rect 224182 693178 224354 693414
rect 223774 693094 224354 693178
rect 223774 692858 223946 693094
rect 224182 692858 224354 693094
rect 223774 657414 224354 692858
rect 223774 657178 223946 657414
rect 224182 657178 224354 657414
rect 223774 657094 224354 657178
rect 223774 656858 223946 657094
rect 224182 656858 224354 657094
rect 223774 621414 224354 656858
rect 223774 621178 223946 621414
rect 224182 621178 224354 621414
rect 223774 621094 224354 621178
rect 223774 620858 223946 621094
rect 224182 620858 224354 621094
rect 223774 585414 224354 620858
rect 223774 585178 223946 585414
rect 224182 585178 224354 585414
rect 223774 585094 224354 585178
rect 223774 584858 223946 585094
rect 224182 584858 224354 585094
rect 223774 549414 224354 584858
rect 223774 549178 223946 549414
rect 224182 549178 224354 549414
rect 223774 549094 224354 549178
rect 223774 548858 223946 549094
rect 224182 548858 224354 549094
rect 223774 513414 224354 548858
rect 223774 513178 223946 513414
rect 224182 513178 224354 513414
rect 223774 513094 224354 513178
rect 223774 512858 223946 513094
rect 224182 512858 224354 513094
rect 223774 477414 224354 512858
rect 223774 477178 223946 477414
rect 224182 477178 224354 477414
rect 223774 477094 224354 477178
rect 223774 476858 223946 477094
rect 224182 476858 224354 477094
rect 223774 441414 224354 476858
rect 223774 441178 223946 441414
rect 224182 441178 224354 441414
rect 223774 441094 224354 441178
rect 223774 440858 223946 441094
rect 224182 440858 224354 441094
rect 223774 405414 224354 440858
rect 223774 405178 223946 405414
rect 224182 405178 224354 405414
rect 223774 405094 224354 405178
rect 223774 404858 223946 405094
rect 224182 404858 224354 405094
rect 223774 369414 224354 404858
rect 223774 369178 223946 369414
rect 224182 369178 224354 369414
rect 223774 369094 224354 369178
rect 223774 368858 223946 369094
rect 224182 368858 224354 369094
rect 223774 333414 224354 368858
rect 223774 333178 223946 333414
rect 224182 333178 224354 333414
rect 223774 333094 224354 333178
rect 223774 332858 223946 333094
rect 224182 332858 224354 333094
rect 223774 297414 224354 332858
rect 223774 297178 223946 297414
rect 224182 297178 224354 297414
rect 223774 297094 224354 297178
rect 223774 296858 223946 297094
rect 224182 296858 224354 297094
rect 223774 261414 224354 296858
rect 223774 261178 223946 261414
rect 224182 261178 224354 261414
rect 223774 261094 224354 261178
rect 223774 260858 223946 261094
rect 224182 260858 224354 261094
rect 223774 225414 224354 260858
rect 223774 225178 223946 225414
rect 224182 225178 224354 225414
rect 223774 225094 224354 225178
rect 223774 224858 223946 225094
rect 224182 224858 224354 225094
rect 223774 189414 224354 224858
rect 223774 189178 223946 189414
rect 224182 189178 224354 189414
rect 223774 189094 224354 189178
rect 223774 188858 223946 189094
rect 224182 188858 224354 189094
rect 223774 153414 224354 188858
rect 223774 153178 223946 153414
rect 224182 153178 224354 153414
rect 223774 153094 224354 153178
rect 223774 152858 223946 153094
rect 224182 152858 224354 153094
rect 223774 117414 224354 152858
rect 223774 117178 223946 117414
rect 224182 117178 224354 117414
rect 223774 117094 224354 117178
rect 223774 116858 223946 117094
rect 224182 116858 224354 117094
rect 223774 81414 224354 116858
rect 223774 81178 223946 81414
rect 224182 81178 224354 81414
rect 223774 81094 224354 81178
rect 223774 80858 223946 81094
rect 224182 80858 224354 81094
rect 223774 45414 224354 80858
rect 223774 45178 223946 45414
rect 224182 45178 224354 45414
rect 223774 45094 224354 45178
rect 223774 44858 223946 45094
rect 224182 44858 224354 45094
rect 223774 9414 224354 44858
rect 223774 9178 223946 9414
rect 224182 9178 224354 9414
rect 223774 9094 224354 9178
rect 223774 8858 223946 9094
rect 224182 8858 224354 9094
rect 223774 -4026 224354 8858
rect 223774 -4262 223946 -4026
rect 224182 -4262 224354 -4026
rect 223774 -4346 224354 -4262
rect 223774 -4582 223946 -4346
rect 224182 -4582 224354 -4346
rect 223774 -5514 224354 -4582
rect 227254 696894 227834 709802
rect 245254 711278 245834 711290
rect 245254 711042 245426 711278
rect 245662 711042 245834 711278
rect 245254 710958 245834 711042
rect 245254 710722 245426 710958
rect 245662 710722 245834 710958
rect 241774 709438 242354 709450
rect 241774 709202 241946 709438
rect 242182 709202 242354 709438
rect 241774 709118 242354 709202
rect 241774 708882 241946 709118
rect 242182 708882 242354 709118
rect 238294 707598 238874 707610
rect 238294 707362 238466 707598
rect 238702 707362 238874 707598
rect 238294 707278 238874 707362
rect 238294 707042 238466 707278
rect 238702 707042 238874 707278
rect 227254 696658 227426 696894
rect 227662 696658 227834 696894
rect 227254 696574 227834 696658
rect 227254 696338 227426 696574
rect 227662 696338 227834 696574
rect 227254 660894 227834 696338
rect 227254 660658 227426 660894
rect 227662 660658 227834 660894
rect 227254 660574 227834 660658
rect 227254 660338 227426 660574
rect 227662 660338 227834 660574
rect 227254 624894 227834 660338
rect 227254 624658 227426 624894
rect 227662 624658 227834 624894
rect 227254 624574 227834 624658
rect 227254 624338 227426 624574
rect 227662 624338 227834 624574
rect 227254 588894 227834 624338
rect 227254 588658 227426 588894
rect 227662 588658 227834 588894
rect 227254 588574 227834 588658
rect 227254 588338 227426 588574
rect 227662 588338 227834 588574
rect 227254 552894 227834 588338
rect 227254 552658 227426 552894
rect 227662 552658 227834 552894
rect 227254 552574 227834 552658
rect 227254 552338 227426 552574
rect 227662 552338 227834 552574
rect 227254 516894 227834 552338
rect 227254 516658 227426 516894
rect 227662 516658 227834 516894
rect 227254 516574 227834 516658
rect 227254 516338 227426 516574
rect 227662 516338 227834 516574
rect 227254 480894 227834 516338
rect 227254 480658 227426 480894
rect 227662 480658 227834 480894
rect 227254 480574 227834 480658
rect 227254 480338 227426 480574
rect 227662 480338 227834 480574
rect 227254 444894 227834 480338
rect 227254 444658 227426 444894
rect 227662 444658 227834 444894
rect 227254 444574 227834 444658
rect 227254 444338 227426 444574
rect 227662 444338 227834 444574
rect 227254 408894 227834 444338
rect 227254 408658 227426 408894
rect 227662 408658 227834 408894
rect 227254 408574 227834 408658
rect 227254 408338 227426 408574
rect 227662 408338 227834 408574
rect 227254 372894 227834 408338
rect 227254 372658 227426 372894
rect 227662 372658 227834 372894
rect 227254 372574 227834 372658
rect 227254 372338 227426 372574
rect 227662 372338 227834 372574
rect 227254 336894 227834 372338
rect 234814 705758 235394 705770
rect 234814 705522 234986 705758
rect 235222 705522 235394 705758
rect 234814 705438 235394 705522
rect 234814 705202 234986 705438
rect 235222 705202 235394 705438
rect 234814 668454 235394 705202
rect 234814 668218 234986 668454
rect 235222 668218 235394 668454
rect 234814 668134 235394 668218
rect 234814 667898 234986 668134
rect 235222 667898 235394 668134
rect 234814 632454 235394 667898
rect 234814 632218 234986 632454
rect 235222 632218 235394 632454
rect 234814 632134 235394 632218
rect 234814 631898 234986 632134
rect 235222 631898 235394 632134
rect 234814 596454 235394 631898
rect 234814 596218 234986 596454
rect 235222 596218 235394 596454
rect 234814 596134 235394 596218
rect 234814 595898 234986 596134
rect 235222 595898 235394 596134
rect 234814 560454 235394 595898
rect 234814 560218 234986 560454
rect 235222 560218 235394 560454
rect 234814 560134 235394 560218
rect 234814 559898 234986 560134
rect 235222 559898 235394 560134
rect 234814 524454 235394 559898
rect 234814 524218 234986 524454
rect 235222 524218 235394 524454
rect 234814 524134 235394 524218
rect 234814 523898 234986 524134
rect 235222 523898 235394 524134
rect 234814 488454 235394 523898
rect 234814 488218 234986 488454
rect 235222 488218 235394 488454
rect 234814 488134 235394 488218
rect 234814 487898 234986 488134
rect 235222 487898 235394 488134
rect 234814 452454 235394 487898
rect 234814 452218 234986 452454
rect 235222 452218 235394 452454
rect 234814 452134 235394 452218
rect 234814 451898 234986 452134
rect 235222 451898 235394 452134
rect 234814 416454 235394 451898
rect 234814 416218 234986 416454
rect 235222 416218 235394 416454
rect 234814 416134 235394 416218
rect 234814 415898 234986 416134
rect 235222 415898 235394 416134
rect 234814 380454 235394 415898
rect 234814 380218 234986 380454
rect 235222 380218 235394 380454
rect 234814 380134 235394 380218
rect 234814 379898 234986 380134
rect 235222 379898 235394 380134
rect 230795 361180 230861 361181
rect 230795 361116 230796 361180
rect 230860 361116 230861 361180
rect 230795 361115 230861 361116
rect 230798 360858 230858 361115
rect 227254 336658 227426 336894
rect 227662 336658 227834 336894
rect 227254 336574 227834 336658
rect 227254 336338 227426 336574
rect 227662 336338 227834 336574
rect 227254 300894 227834 336338
rect 227254 300658 227426 300894
rect 227662 300658 227834 300894
rect 227254 300574 227834 300658
rect 227254 300338 227426 300574
rect 227662 300338 227834 300574
rect 227254 264894 227834 300338
rect 227254 264658 227426 264894
rect 227662 264658 227834 264894
rect 227254 264574 227834 264658
rect 227254 264338 227426 264574
rect 227662 264338 227834 264574
rect 227254 228894 227834 264338
rect 227254 228658 227426 228894
rect 227662 228658 227834 228894
rect 227254 228574 227834 228658
rect 227254 228338 227426 228574
rect 227662 228338 227834 228574
rect 227254 192894 227834 228338
rect 227254 192658 227426 192894
rect 227662 192658 227834 192894
rect 227254 192574 227834 192658
rect 227254 192338 227426 192574
rect 227662 192338 227834 192574
rect 227254 156894 227834 192338
rect 227254 156658 227426 156894
rect 227662 156658 227834 156894
rect 227254 156574 227834 156658
rect 227254 156338 227426 156574
rect 227662 156338 227834 156574
rect 227254 120894 227834 156338
rect 227254 120658 227426 120894
rect 227662 120658 227834 120894
rect 227254 120574 227834 120658
rect 227254 120338 227426 120574
rect 227662 120338 227834 120574
rect 227254 84894 227834 120338
rect 227254 84658 227426 84894
rect 227662 84658 227834 84894
rect 227254 84574 227834 84658
rect 227254 84338 227426 84574
rect 227662 84338 227834 84574
rect 227254 48894 227834 84338
rect 227254 48658 227426 48894
rect 227662 48658 227834 48894
rect 227254 48574 227834 48658
rect 227254 48338 227426 48574
rect 227662 48338 227834 48574
rect 227254 12894 227834 48338
rect 227254 12658 227426 12894
rect 227662 12658 227834 12894
rect 227254 12574 227834 12658
rect 227254 12338 227426 12574
rect 227662 12338 227834 12574
rect 209254 -7022 209426 -6786
rect 209662 -7022 209834 -6786
rect 209254 -7106 209834 -7022
rect 209254 -7342 209426 -7106
rect 209662 -7342 209834 -7106
rect 209254 -7354 209834 -7342
rect 227254 -5866 227834 12338
rect 234814 344454 235394 379898
rect 234814 344218 234986 344454
rect 235222 344218 235394 344454
rect 234814 344134 235394 344218
rect 234814 343898 234986 344134
rect 235222 343898 235394 344134
rect 234814 308454 235394 343898
rect 234814 308218 234986 308454
rect 235222 308218 235394 308454
rect 234814 308134 235394 308218
rect 234814 307898 234986 308134
rect 235222 307898 235394 308134
rect 234814 272454 235394 307898
rect 234814 272218 234986 272454
rect 235222 272218 235394 272454
rect 234814 272134 235394 272218
rect 234814 271898 234986 272134
rect 235222 271898 235394 272134
rect 234814 236454 235394 271898
rect 234814 236218 234986 236454
rect 235222 236218 235394 236454
rect 234814 236134 235394 236218
rect 234814 235898 234986 236134
rect 235222 235898 235394 236134
rect 234814 200454 235394 235898
rect 234814 200218 234986 200454
rect 235222 200218 235394 200454
rect 234814 200134 235394 200218
rect 234814 199898 234986 200134
rect 235222 199898 235394 200134
rect 234814 164454 235394 199898
rect 234814 164218 234986 164454
rect 235222 164218 235394 164454
rect 234814 164134 235394 164218
rect 234814 163898 234986 164134
rect 235222 163898 235394 164134
rect 234814 128454 235394 163898
rect 234814 128218 234986 128454
rect 235222 128218 235394 128454
rect 234814 128134 235394 128218
rect 234814 127898 234986 128134
rect 235222 127898 235394 128134
rect 234814 92454 235394 127898
rect 234814 92218 234986 92454
rect 235222 92218 235394 92454
rect 234814 92134 235394 92218
rect 234814 91898 234986 92134
rect 235222 91898 235394 92134
rect 234814 56454 235394 91898
rect 234814 56218 234986 56454
rect 235222 56218 235394 56454
rect 234814 56134 235394 56218
rect 234814 55898 234986 56134
rect 235222 55898 235394 56134
rect 234814 20454 235394 55898
rect 234814 20218 234986 20454
rect 235222 20218 235394 20454
rect 234814 20134 235394 20218
rect 234814 19898 234986 20134
rect 235222 19898 235394 20134
rect 234814 -1266 235394 19898
rect 234814 -1502 234986 -1266
rect 235222 -1502 235394 -1266
rect 234814 -1586 235394 -1502
rect 234814 -1822 234986 -1586
rect 235222 -1822 235394 -1586
rect 234814 -1834 235394 -1822
rect 238294 671934 238874 707042
rect 238294 671698 238466 671934
rect 238702 671698 238874 671934
rect 238294 671614 238874 671698
rect 238294 671378 238466 671614
rect 238702 671378 238874 671614
rect 238294 635934 238874 671378
rect 238294 635698 238466 635934
rect 238702 635698 238874 635934
rect 238294 635614 238874 635698
rect 238294 635378 238466 635614
rect 238702 635378 238874 635614
rect 238294 599934 238874 635378
rect 238294 599698 238466 599934
rect 238702 599698 238874 599934
rect 238294 599614 238874 599698
rect 238294 599378 238466 599614
rect 238702 599378 238874 599614
rect 238294 563934 238874 599378
rect 238294 563698 238466 563934
rect 238702 563698 238874 563934
rect 238294 563614 238874 563698
rect 238294 563378 238466 563614
rect 238702 563378 238874 563614
rect 238294 527934 238874 563378
rect 238294 527698 238466 527934
rect 238702 527698 238874 527934
rect 238294 527614 238874 527698
rect 238294 527378 238466 527614
rect 238702 527378 238874 527614
rect 238294 491934 238874 527378
rect 238294 491698 238466 491934
rect 238702 491698 238874 491934
rect 238294 491614 238874 491698
rect 238294 491378 238466 491614
rect 238702 491378 238874 491614
rect 238294 455934 238874 491378
rect 238294 455698 238466 455934
rect 238702 455698 238874 455934
rect 238294 455614 238874 455698
rect 238294 455378 238466 455614
rect 238702 455378 238874 455614
rect 238294 419934 238874 455378
rect 238294 419698 238466 419934
rect 238702 419698 238874 419934
rect 238294 419614 238874 419698
rect 238294 419378 238466 419614
rect 238702 419378 238874 419614
rect 238294 383934 238874 419378
rect 238294 383698 238466 383934
rect 238702 383698 238874 383934
rect 238294 383614 238874 383698
rect 238294 383378 238466 383614
rect 238702 383378 238874 383614
rect 238294 347934 238874 383378
rect 241774 675414 242354 708882
rect 241774 675178 241946 675414
rect 242182 675178 242354 675414
rect 241774 675094 242354 675178
rect 241774 674858 241946 675094
rect 242182 674858 242354 675094
rect 241774 639414 242354 674858
rect 241774 639178 241946 639414
rect 242182 639178 242354 639414
rect 241774 639094 242354 639178
rect 241774 638858 241946 639094
rect 242182 638858 242354 639094
rect 241774 603414 242354 638858
rect 241774 603178 241946 603414
rect 242182 603178 242354 603414
rect 241774 603094 242354 603178
rect 241774 602858 241946 603094
rect 242182 602858 242354 603094
rect 241774 567414 242354 602858
rect 241774 567178 241946 567414
rect 242182 567178 242354 567414
rect 241774 567094 242354 567178
rect 241774 566858 241946 567094
rect 242182 566858 242354 567094
rect 241774 531414 242354 566858
rect 241774 531178 241946 531414
rect 242182 531178 242354 531414
rect 241774 531094 242354 531178
rect 241774 530858 241946 531094
rect 242182 530858 242354 531094
rect 241774 495414 242354 530858
rect 241774 495178 241946 495414
rect 242182 495178 242354 495414
rect 241774 495094 242354 495178
rect 241774 494858 241946 495094
rect 242182 494858 242354 495094
rect 241774 459414 242354 494858
rect 241774 459178 241946 459414
rect 242182 459178 242354 459414
rect 241774 459094 242354 459178
rect 241774 458858 241946 459094
rect 242182 458858 242354 459094
rect 241774 423414 242354 458858
rect 241774 423178 241946 423414
rect 242182 423178 242354 423414
rect 241774 423094 242354 423178
rect 241774 422858 241946 423094
rect 242182 422858 242354 423094
rect 241774 387414 242354 422858
rect 241774 387178 241946 387414
rect 242182 387178 242354 387414
rect 241774 387094 242354 387178
rect 241774 386858 241946 387094
rect 242182 386858 242354 387094
rect 239078 360858 239138 363342
rect 238294 347698 238466 347934
rect 238702 347698 238874 347934
rect 238294 347614 238874 347698
rect 238294 347378 238466 347614
rect 238702 347378 238874 347614
rect 238294 311934 238874 347378
rect 238294 311698 238466 311934
rect 238702 311698 238874 311934
rect 238294 311614 238874 311698
rect 238294 311378 238466 311614
rect 238702 311378 238874 311614
rect 238294 275934 238874 311378
rect 238294 275698 238466 275934
rect 238702 275698 238874 275934
rect 238294 275614 238874 275698
rect 238294 275378 238466 275614
rect 238702 275378 238874 275614
rect 238294 239934 238874 275378
rect 238294 239698 238466 239934
rect 238702 239698 238874 239934
rect 238294 239614 238874 239698
rect 238294 239378 238466 239614
rect 238702 239378 238874 239614
rect 238294 203934 238874 239378
rect 238294 203698 238466 203934
rect 238702 203698 238874 203934
rect 238294 203614 238874 203698
rect 238294 203378 238466 203614
rect 238702 203378 238874 203614
rect 238294 167934 238874 203378
rect 238294 167698 238466 167934
rect 238702 167698 238874 167934
rect 238294 167614 238874 167698
rect 238294 167378 238466 167614
rect 238702 167378 238874 167614
rect 238294 131934 238874 167378
rect 238294 131698 238466 131934
rect 238702 131698 238874 131934
rect 238294 131614 238874 131698
rect 238294 131378 238466 131614
rect 238702 131378 238874 131614
rect 238294 95934 238874 131378
rect 238294 95698 238466 95934
rect 238702 95698 238874 95934
rect 238294 95614 238874 95698
rect 238294 95378 238466 95614
rect 238702 95378 238874 95614
rect 238294 59934 238874 95378
rect 238294 59698 238466 59934
rect 238702 59698 238874 59934
rect 238294 59614 238874 59698
rect 238294 59378 238466 59614
rect 238702 59378 238874 59614
rect 238294 23934 238874 59378
rect 238294 23698 238466 23934
rect 238702 23698 238874 23934
rect 238294 23614 238874 23698
rect 238294 23378 238466 23614
rect 238702 23378 238874 23614
rect 238294 -3106 238874 23378
rect 238294 -3342 238466 -3106
rect 238702 -3342 238874 -3106
rect 238294 -3426 238874 -3342
rect 238294 -3662 238466 -3426
rect 238702 -3662 238874 -3426
rect 238294 -3674 238874 -3662
rect 241774 351414 242354 386858
rect 241774 351178 241946 351414
rect 242182 351178 242354 351414
rect 241774 351094 242354 351178
rect 241774 350858 241946 351094
rect 242182 350858 242354 351094
rect 241774 315414 242354 350858
rect 241774 315178 241946 315414
rect 242182 315178 242354 315414
rect 241774 315094 242354 315178
rect 241774 314858 241946 315094
rect 242182 314858 242354 315094
rect 241774 279414 242354 314858
rect 241774 279178 241946 279414
rect 242182 279178 242354 279414
rect 241774 279094 242354 279178
rect 241774 278858 241946 279094
rect 242182 278858 242354 279094
rect 241774 243414 242354 278858
rect 241774 243178 241946 243414
rect 242182 243178 242354 243414
rect 241774 243094 242354 243178
rect 241774 242858 241946 243094
rect 242182 242858 242354 243094
rect 241774 207414 242354 242858
rect 241774 207178 241946 207414
rect 242182 207178 242354 207414
rect 241774 207094 242354 207178
rect 241774 206858 241946 207094
rect 242182 206858 242354 207094
rect 241774 171414 242354 206858
rect 241774 171178 241946 171414
rect 242182 171178 242354 171414
rect 241774 171094 242354 171178
rect 241774 170858 241946 171094
rect 242182 170858 242354 171094
rect 241774 135414 242354 170858
rect 241774 135178 241946 135414
rect 242182 135178 242354 135414
rect 241774 135094 242354 135178
rect 241774 134858 241946 135094
rect 242182 134858 242354 135094
rect 241774 99414 242354 134858
rect 241774 99178 241946 99414
rect 242182 99178 242354 99414
rect 241774 99094 242354 99178
rect 241774 98858 241946 99094
rect 242182 98858 242354 99094
rect 241774 63414 242354 98858
rect 241774 63178 241946 63414
rect 242182 63178 242354 63414
rect 241774 63094 242354 63178
rect 241774 62858 241946 63094
rect 242182 62858 242354 63094
rect 241774 27414 242354 62858
rect 241774 27178 241946 27414
rect 242182 27178 242354 27414
rect 241774 27094 242354 27178
rect 241774 26858 241946 27094
rect 242182 26858 242354 27094
rect 241774 -4946 242354 26858
rect 241774 -5182 241946 -4946
rect 242182 -5182 242354 -4946
rect 241774 -5266 242354 -5182
rect 241774 -5502 241946 -5266
rect 242182 -5502 242354 -5266
rect 241774 -5514 242354 -5502
rect 245254 678894 245834 710722
rect 263254 710358 263834 711290
rect 263254 710122 263426 710358
rect 263662 710122 263834 710358
rect 263254 710038 263834 710122
rect 263254 709802 263426 710038
rect 263662 709802 263834 710038
rect 259774 708518 260354 709450
rect 259774 708282 259946 708518
rect 260182 708282 260354 708518
rect 259774 708198 260354 708282
rect 259774 707962 259946 708198
rect 260182 707962 260354 708198
rect 256294 706678 256874 707610
rect 256294 706442 256466 706678
rect 256702 706442 256874 706678
rect 256294 706358 256874 706442
rect 256294 706122 256466 706358
rect 256702 706122 256874 706358
rect 245254 678658 245426 678894
rect 245662 678658 245834 678894
rect 245254 678574 245834 678658
rect 245254 678338 245426 678574
rect 245662 678338 245834 678574
rect 245254 642894 245834 678338
rect 245254 642658 245426 642894
rect 245662 642658 245834 642894
rect 245254 642574 245834 642658
rect 245254 642338 245426 642574
rect 245662 642338 245834 642574
rect 245254 606894 245834 642338
rect 245254 606658 245426 606894
rect 245662 606658 245834 606894
rect 245254 606574 245834 606658
rect 245254 606338 245426 606574
rect 245662 606338 245834 606574
rect 245254 570894 245834 606338
rect 245254 570658 245426 570894
rect 245662 570658 245834 570894
rect 245254 570574 245834 570658
rect 245254 570338 245426 570574
rect 245662 570338 245834 570574
rect 245254 534894 245834 570338
rect 245254 534658 245426 534894
rect 245662 534658 245834 534894
rect 245254 534574 245834 534658
rect 245254 534338 245426 534574
rect 245662 534338 245834 534574
rect 245254 498894 245834 534338
rect 245254 498658 245426 498894
rect 245662 498658 245834 498894
rect 245254 498574 245834 498658
rect 245254 498338 245426 498574
rect 245662 498338 245834 498574
rect 245254 462894 245834 498338
rect 245254 462658 245426 462894
rect 245662 462658 245834 462894
rect 245254 462574 245834 462658
rect 245254 462338 245426 462574
rect 245662 462338 245834 462574
rect 245254 426894 245834 462338
rect 245254 426658 245426 426894
rect 245662 426658 245834 426894
rect 245254 426574 245834 426658
rect 245254 426338 245426 426574
rect 245662 426338 245834 426574
rect 245254 390894 245834 426338
rect 245254 390658 245426 390894
rect 245662 390658 245834 390894
rect 245254 390574 245834 390658
rect 245254 390338 245426 390574
rect 245662 390338 245834 390574
rect 245254 354894 245834 390338
rect 252814 704838 253394 705770
rect 252814 704602 252986 704838
rect 253222 704602 253394 704838
rect 252814 704518 253394 704602
rect 252814 704282 252986 704518
rect 253222 704282 253394 704518
rect 252814 686454 253394 704282
rect 252814 686218 252986 686454
rect 253222 686218 253394 686454
rect 252814 686134 253394 686218
rect 252814 685898 252986 686134
rect 253222 685898 253394 686134
rect 252814 650454 253394 685898
rect 252814 650218 252986 650454
rect 253222 650218 253394 650454
rect 252814 650134 253394 650218
rect 252814 649898 252986 650134
rect 253222 649898 253394 650134
rect 252814 614454 253394 649898
rect 252814 614218 252986 614454
rect 253222 614218 253394 614454
rect 252814 614134 253394 614218
rect 252814 613898 252986 614134
rect 253222 613898 253394 614134
rect 252814 578454 253394 613898
rect 252814 578218 252986 578454
rect 253222 578218 253394 578454
rect 252814 578134 253394 578218
rect 252814 577898 252986 578134
rect 253222 577898 253394 578134
rect 252814 542454 253394 577898
rect 252814 542218 252986 542454
rect 253222 542218 253394 542454
rect 252814 542134 253394 542218
rect 252814 541898 252986 542134
rect 253222 541898 253394 542134
rect 252814 506454 253394 541898
rect 252814 506218 252986 506454
rect 253222 506218 253394 506454
rect 252814 506134 253394 506218
rect 252814 505898 252986 506134
rect 253222 505898 253394 506134
rect 252814 470454 253394 505898
rect 252814 470218 252986 470454
rect 253222 470218 253394 470454
rect 252814 470134 253394 470218
rect 252814 469898 252986 470134
rect 253222 469898 253394 470134
rect 252814 434454 253394 469898
rect 252814 434218 252986 434454
rect 253222 434218 253394 434454
rect 252814 434134 253394 434218
rect 252814 433898 252986 434134
rect 253222 433898 253394 434134
rect 252814 398454 253394 433898
rect 252814 398218 252986 398454
rect 253222 398218 253394 398454
rect 252814 398134 253394 398218
rect 252814 397898 252986 398134
rect 253222 397898 253394 398134
rect 248646 360858 248706 363342
rect 252814 362454 253394 397898
rect 252814 362218 252986 362454
rect 253222 362218 253394 362454
rect 252814 362134 253394 362218
rect 252814 361898 252986 362134
rect 253222 361898 253394 362134
rect 245254 354658 245426 354894
rect 245662 354658 245834 354894
rect 245254 354574 245834 354658
rect 245254 354338 245426 354574
rect 245662 354338 245834 354574
rect 245254 318894 245834 354338
rect 245254 318658 245426 318894
rect 245662 318658 245834 318894
rect 245254 318574 245834 318658
rect 245254 318338 245426 318574
rect 245662 318338 245834 318574
rect 245254 282894 245834 318338
rect 245254 282658 245426 282894
rect 245662 282658 245834 282894
rect 245254 282574 245834 282658
rect 245254 282338 245426 282574
rect 245662 282338 245834 282574
rect 245254 246894 245834 282338
rect 245254 246658 245426 246894
rect 245662 246658 245834 246894
rect 245254 246574 245834 246658
rect 245254 246338 245426 246574
rect 245662 246338 245834 246574
rect 245254 210894 245834 246338
rect 245254 210658 245426 210894
rect 245662 210658 245834 210894
rect 245254 210574 245834 210658
rect 245254 210338 245426 210574
rect 245662 210338 245834 210574
rect 245254 174894 245834 210338
rect 245254 174658 245426 174894
rect 245662 174658 245834 174894
rect 245254 174574 245834 174658
rect 245254 174338 245426 174574
rect 245662 174338 245834 174574
rect 245254 138894 245834 174338
rect 245254 138658 245426 138894
rect 245662 138658 245834 138894
rect 245254 138574 245834 138658
rect 245254 138338 245426 138574
rect 245662 138338 245834 138574
rect 245254 102894 245834 138338
rect 245254 102658 245426 102894
rect 245662 102658 245834 102894
rect 245254 102574 245834 102658
rect 245254 102338 245426 102574
rect 245662 102338 245834 102574
rect 245254 66894 245834 102338
rect 245254 66658 245426 66894
rect 245662 66658 245834 66894
rect 245254 66574 245834 66658
rect 245254 66338 245426 66574
rect 245662 66338 245834 66574
rect 245254 30894 245834 66338
rect 245254 30658 245426 30894
rect 245662 30658 245834 30894
rect 245254 30574 245834 30658
rect 245254 30338 245426 30574
rect 245662 30338 245834 30574
rect 227254 -6102 227426 -5866
rect 227662 -6102 227834 -5866
rect 227254 -6186 227834 -6102
rect 227254 -6422 227426 -6186
rect 227662 -6422 227834 -6186
rect 227254 -7354 227834 -6422
rect 245254 -6786 245834 30338
rect 252814 326454 253394 361898
rect 252814 326218 252986 326454
rect 253222 326218 253394 326454
rect 252814 326134 253394 326218
rect 252814 325898 252986 326134
rect 253222 325898 253394 326134
rect 252814 290454 253394 325898
rect 252814 290218 252986 290454
rect 253222 290218 253394 290454
rect 252814 290134 253394 290218
rect 252814 289898 252986 290134
rect 253222 289898 253394 290134
rect 252814 254454 253394 289898
rect 252814 254218 252986 254454
rect 253222 254218 253394 254454
rect 252814 254134 253394 254218
rect 252814 253898 252986 254134
rect 253222 253898 253394 254134
rect 252814 218454 253394 253898
rect 252814 218218 252986 218454
rect 253222 218218 253394 218454
rect 252814 218134 253394 218218
rect 252814 217898 252986 218134
rect 253222 217898 253394 218134
rect 252814 182454 253394 217898
rect 252814 182218 252986 182454
rect 253222 182218 253394 182454
rect 252814 182134 253394 182218
rect 252814 181898 252986 182134
rect 253222 181898 253394 182134
rect 252814 146454 253394 181898
rect 252814 146218 252986 146454
rect 253222 146218 253394 146454
rect 252814 146134 253394 146218
rect 252814 145898 252986 146134
rect 253222 145898 253394 146134
rect 252814 110454 253394 145898
rect 252814 110218 252986 110454
rect 253222 110218 253394 110454
rect 252814 110134 253394 110218
rect 252814 109898 252986 110134
rect 253222 109898 253394 110134
rect 252814 74454 253394 109898
rect 252814 74218 252986 74454
rect 253222 74218 253394 74454
rect 252814 74134 253394 74218
rect 252814 73898 252986 74134
rect 253222 73898 253394 74134
rect 252814 38454 253394 73898
rect 252814 38218 252986 38454
rect 253222 38218 253394 38454
rect 252814 38134 253394 38218
rect 252814 37898 252986 38134
rect 253222 37898 253394 38134
rect 252814 2454 253394 37898
rect 252814 2218 252986 2454
rect 253222 2218 253394 2454
rect 252814 2134 253394 2218
rect 252814 1898 252986 2134
rect 253222 1898 253394 2134
rect 252814 -346 253394 1898
rect 252814 -582 252986 -346
rect 253222 -582 253394 -346
rect 252814 -666 253394 -582
rect 252814 -902 252986 -666
rect 253222 -902 253394 -666
rect 252814 -1834 253394 -902
rect 256294 689934 256874 706122
rect 256294 689698 256466 689934
rect 256702 689698 256874 689934
rect 256294 689614 256874 689698
rect 256294 689378 256466 689614
rect 256702 689378 256874 689614
rect 256294 653934 256874 689378
rect 256294 653698 256466 653934
rect 256702 653698 256874 653934
rect 256294 653614 256874 653698
rect 256294 653378 256466 653614
rect 256702 653378 256874 653614
rect 256294 617934 256874 653378
rect 256294 617698 256466 617934
rect 256702 617698 256874 617934
rect 256294 617614 256874 617698
rect 256294 617378 256466 617614
rect 256702 617378 256874 617614
rect 256294 581934 256874 617378
rect 256294 581698 256466 581934
rect 256702 581698 256874 581934
rect 256294 581614 256874 581698
rect 256294 581378 256466 581614
rect 256702 581378 256874 581614
rect 256294 545934 256874 581378
rect 256294 545698 256466 545934
rect 256702 545698 256874 545934
rect 256294 545614 256874 545698
rect 256294 545378 256466 545614
rect 256702 545378 256874 545614
rect 256294 509934 256874 545378
rect 256294 509698 256466 509934
rect 256702 509698 256874 509934
rect 256294 509614 256874 509698
rect 256294 509378 256466 509614
rect 256702 509378 256874 509614
rect 256294 473934 256874 509378
rect 256294 473698 256466 473934
rect 256702 473698 256874 473934
rect 256294 473614 256874 473698
rect 256294 473378 256466 473614
rect 256702 473378 256874 473614
rect 256294 437934 256874 473378
rect 256294 437698 256466 437934
rect 256702 437698 256874 437934
rect 256294 437614 256874 437698
rect 256294 437378 256466 437614
rect 256702 437378 256874 437614
rect 256294 401934 256874 437378
rect 256294 401698 256466 401934
rect 256702 401698 256874 401934
rect 256294 401614 256874 401698
rect 256294 401378 256466 401614
rect 256702 401378 256874 401614
rect 256294 365934 256874 401378
rect 256294 365698 256466 365934
rect 256702 365698 256874 365934
rect 256294 365614 256874 365698
rect 256294 365378 256466 365614
rect 256702 365378 256874 365614
rect 256294 329934 256874 365378
rect 256294 329698 256466 329934
rect 256702 329698 256874 329934
rect 256294 329614 256874 329698
rect 256294 329378 256466 329614
rect 256702 329378 256874 329614
rect 256294 293934 256874 329378
rect 256294 293698 256466 293934
rect 256702 293698 256874 293934
rect 256294 293614 256874 293698
rect 256294 293378 256466 293614
rect 256702 293378 256874 293614
rect 256294 257934 256874 293378
rect 256294 257698 256466 257934
rect 256702 257698 256874 257934
rect 256294 257614 256874 257698
rect 256294 257378 256466 257614
rect 256702 257378 256874 257614
rect 256294 221934 256874 257378
rect 256294 221698 256466 221934
rect 256702 221698 256874 221934
rect 256294 221614 256874 221698
rect 256294 221378 256466 221614
rect 256702 221378 256874 221614
rect 256294 185934 256874 221378
rect 256294 185698 256466 185934
rect 256702 185698 256874 185934
rect 256294 185614 256874 185698
rect 256294 185378 256466 185614
rect 256702 185378 256874 185614
rect 256294 149934 256874 185378
rect 256294 149698 256466 149934
rect 256702 149698 256874 149934
rect 256294 149614 256874 149698
rect 256294 149378 256466 149614
rect 256702 149378 256874 149614
rect 256294 113934 256874 149378
rect 256294 113698 256466 113934
rect 256702 113698 256874 113934
rect 256294 113614 256874 113698
rect 256294 113378 256466 113614
rect 256702 113378 256874 113614
rect 256294 77934 256874 113378
rect 256294 77698 256466 77934
rect 256702 77698 256874 77934
rect 256294 77614 256874 77698
rect 256294 77378 256466 77614
rect 256702 77378 256874 77614
rect 256294 41934 256874 77378
rect 256294 41698 256466 41934
rect 256702 41698 256874 41934
rect 256294 41614 256874 41698
rect 256294 41378 256466 41614
rect 256702 41378 256874 41614
rect 256294 5934 256874 41378
rect 256294 5698 256466 5934
rect 256702 5698 256874 5934
rect 256294 5614 256874 5698
rect 256294 5378 256466 5614
rect 256702 5378 256874 5614
rect 256294 -2186 256874 5378
rect 256294 -2422 256466 -2186
rect 256702 -2422 256874 -2186
rect 256294 -2506 256874 -2422
rect 256294 -2742 256466 -2506
rect 256702 -2742 256874 -2506
rect 256294 -3674 256874 -2742
rect 259774 693414 260354 707962
rect 259774 693178 259946 693414
rect 260182 693178 260354 693414
rect 259774 693094 260354 693178
rect 259774 692858 259946 693094
rect 260182 692858 260354 693094
rect 259774 657414 260354 692858
rect 259774 657178 259946 657414
rect 260182 657178 260354 657414
rect 259774 657094 260354 657178
rect 259774 656858 259946 657094
rect 260182 656858 260354 657094
rect 259774 621414 260354 656858
rect 259774 621178 259946 621414
rect 260182 621178 260354 621414
rect 259774 621094 260354 621178
rect 259774 620858 259946 621094
rect 260182 620858 260354 621094
rect 259774 585414 260354 620858
rect 259774 585178 259946 585414
rect 260182 585178 260354 585414
rect 259774 585094 260354 585178
rect 259774 584858 259946 585094
rect 260182 584858 260354 585094
rect 259774 549414 260354 584858
rect 259774 549178 259946 549414
rect 260182 549178 260354 549414
rect 259774 549094 260354 549178
rect 259774 548858 259946 549094
rect 260182 548858 260354 549094
rect 259774 513414 260354 548858
rect 259774 513178 259946 513414
rect 260182 513178 260354 513414
rect 259774 513094 260354 513178
rect 259774 512858 259946 513094
rect 260182 512858 260354 513094
rect 259774 477414 260354 512858
rect 259774 477178 259946 477414
rect 260182 477178 260354 477414
rect 259774 477094 260354 477178
rect 259774 476858 259946 477094
rect 260182 476858 260354 477094
rect 259774 441414 260354 476858
rect 259774 441178 259946 441414
rect 260182 441178 260354 441414
rect 259774 441094 260354 441178
rect 259774 440858 259946 441094
rect 260182 440858 260354 441094
rect 259774 405414 260354 440858
rect 259774 405178 259946 405414
rect 260182 405178 260354 405414
rect 259774 405094 260354 405178
rect 259774 404858 259946 405094
rect 260182 404858 260354 405094
rect 259774 369414 260354 404858
rect 259774 369178 259946 369414
rect 260182 369178 260354 369414
rect 259774 369094 260354 369178
rect 259774 368858 259946 369094
rect 260182 368858 260354 369094
rect 259774 333414 260354 368858
rect 259774 333178 259946 333414
rect 260182 333178 260354 333414
rect 259774 333094 260354 333178
rect 259774 332858 259946 333094
rect 260182 332858 260354 333094
rect 259774 297414 260354 332858
rect 259774 297178 259946 297414
rect 260182 297178 260354 297414
rect 259774 297094 260354 297178
rect 259774 296858 259946 297094
rect 260182 296858 260354 297094
rect 259774 261414 260354 296858
rect 259774 261178 259946 261414
rect 260182 261178 260354 261414
rect 259774 261094 260354 261178
rect 259774 260858 259946 261094
rect 260182 260858 260354 261094
rect 259774 225414 260354 260858
rect 259774 225178 259946 225414
rect 260182 225178 260354 225414
rect 259774 225094 260354 225178
rect 259774 224858 259946 225094
rect 260182 224858 260354 225094
rect 259774 189414 260354 224858
rect 259774 189178 259946 189414
rect 260182 189178 260354 189414
rect 259774 189094 260354 189178
rect 259774 188858 259946 189094
rect 260182 188858 260354 189094
rect 259774 153414 260354 188858
rect 259774 153178 259946 153414
rect 260182 153178 260354 153414
rect 259774 153094 260354 153178
rect 259774 152858 259946 153094
rect 260182 152858 260354 153094
rect 259774 117414 260354 152858
rect 259774 117178 259946 117414
rect 260182 117178 260354 117414
rect 259774 117094 260354 117178
rect 259774 116858 259946 117094
rect 260182 116858 260354 117094
rect 259774 81414 260354 116858
rect 259774 81178 259946 81414
rect 260182 81178 260354 81414
rect 259774 81094 260354 81178
rect 259774 80858 259946 81094
rect 260182 80858 260354 81094
rect 259774 45414 260354 80858
rect 259774 45178 259946 45414
rect 260182 45178 260354 45414
rect 259774 45094 260354 45178
rect 259774 44858 259946 45094
rect 260182 44858 260354 45094
rect 259774 9414 260354 44858
rect 259774 9178 259946 9414
rect 260182 9178 260354 9414
rect 259774 9094 260354 9178
rect 259774 8858 259946 9094
rect 260182 8858 260354 9094
rect 259774 -4026 260354 8858
rect 259774 -4262 259946 -4026
rect 260182 -4262 260354 -4026
rect 259774 -4346 260354 -4262
rect 259774 -4582 259946 -4346
rect 260182 -4582 260354 -4346
rect 259774 -5514 260354 -4582
rect 263254 696894 263834 709802
rect 281254 711278 281834 711290
rect 281254 711042 281426 711278
rect 281662 711042 281834 711278
rect 281254 710958 281834 711042
rect 281254 710722 281426 710958
rect 281662 710722 281834 710958
rect 277774 709438 278354 709450
rect 277774 709202 277946 709438
rect 278182 709202 278354 709438
rect 277774 709118 278354 709202
rect 277774 708882 277946 709118
rect 278182 708882 278354 709118
rect 274294 707598 274874 707610
rect 274294 707362 274466 707598
rect 274702 707362 274874 707598
rect 274294 707278 274874 707362
rect 274294 707042 274466 707278
rect 274702 707042 274874 707278
rect 263254 696658 263426 696894
rect 263662 696658 263834 696894
rect 263254 696574 263834 696658
rect 263254 696338 263426 696574
rect 263662 696338 263834 696574
rect 263254 660894 263834 696338
rect 263254 660658 263426 660894
rect 263662 660658 263834 660894
rect 263254 660574 263834 660658
rect 263254 660338 263426 660574
rect 263662 660338 263834 660574
rect 263254 624894 263834 660338
rect 263254 624658 263426 624894
rect 263662 624658 263834 624894
rect 263254 624574 263834 624658
rect 263254 624338 263426 624574
rect 263662 624338 263834 624574
rect 263254 588894 263834 624338
rect 263254 588658 263426 588894
rect 263662 588658 263834 588894
rect 263254 588574 263834 588658
rect 263254 588338 263426 588574
rect 263662 588338 263834 588574
rect 263254 552894 263834 588338
rect 263254 552658 263426 552894
rect 263662 552658 263834 552894
rect 263254 552574 263834 552658
rect 263254 552338 263426 552574
rect 263662 552338 263834 552574
rect 263254 516894 263834 552338
rect 263254 516658 263426 516894
rect 263662 516658 263834 516894
rect 263254 516574 263834 516658
rect 263254 516338 263426 516574
rect 263662 516338 263834 516574
rect 263254 480894 263834 516338
rect 263254 480658 263426 480894
rect 263662 480658 263834 480894
rect 263254 480574 263834 480658
rect 263254 480338 263426 480574
rect 263662 480338 263834 480574
rect 263254 444894 263834 480338
rect 270814 705758 271394 705770
rect 270814 705522 270986 705758
rect 271222 705522 271394 705758
rect 270814 705438 271394 705522
rect 270814 705202 270986 705438
rect 271222 705202 271394 705438
rect 270814 668454 271394 705202
rect 270814 668218 270986 668454
rect 271222 668218 271394 668454
rect 270814 668134 271394 668218
rect 270814 667898 270986 668134
rect 271222 667898 271394 668134
rect 270814 632454 271394 667898
rect 270814 632218 270986 632454
rect 271222 632218 271394 632454
rect 270814 632134 271394 632218
rect 270814 631898 270986 632134
rect 271222 631898 271394 632134
rect 270814 596454 271394 631898
rect 270814 596218 270986 596454
rect 271222 596218 271394 596454
rect 270814 596134 271394 596218
rect 270814 595898 270986 596134
rect 271222 595898 271394 596134
rect 270814 560454 271394 595898
rect 270814 560218 270986 560454
rect 271222 560218 271394 560454
rect 270814 560134 271394 560218
rect 270814 559898 270986 560134
rect 271222 559898 271394 560134
rect 270814 524454 271394 559898
rect 270814 524218 270986 524454
rect 271222 524218 271394 524454
rect 270814 524134 271394 524218
rect 270814 523898 270986 524134
rect 271222 523898 271394 524134
rect 270814 488454 271394 523898
rect 270814 488218 270986 488454
rect 271222 488218 271394 488454
rect 270814 488134 271394 488218
rect 270814 487898 270986 488134
rect 271222 487898 271394 488134
rect 268331 472020 268397 472021
rect 268331 471956 268332 472020
rect 268396 471956 268397 472020
rect 268331 471955 268397 471956
rect 263254 444658 263426 444894
rect 263662 444658 263834 444894
rect 263254 444574 263834 444658
rect 263254 444338 263426 444574
rect 263662 444338 263834 444574
rect 263254 408894 263834 444338
rect 263254 408658 263426 408894
rect 263662 408658 263834 408894
rect 263254 408574 263834 408658
rect 263254 408338 263426 408574
rect 263662 408338 263834 408574
rect 263254 372894 263834 408338
rect 263254 372658 263426 372894
rect 263662 372658 263834 372894
rect 263254 372574 263834 372658
rect 263254 372338 263426 372574
rect 263662 372338 263834 372574
rect 263254 336894 263834 372338
rect 263254 336658 263426 336894
rect 263662 336658 263834 336894
rect 263254 336574 263834 336658
rect 263254 336338 263426 336574
rect 263662 336338 263834 336574
rect 263254 300894 263834 336338
rect 263254 300658 263426 300894
rect 263662 300658 263834 300894
rect 263254 300574 263834 300658
rect 263254 300338 263426 300574
rect 263662 300338 263834 300574
rect 263254 264894 263834 300338
rect 263254 264658 263426 264894
rect 263662 264658 263834 264894
rect 263254 264574 263834 264658
rect 263254 264338 263426 264574
rect 263662 264338 263834 264574
rect 263254 228894 263834 264338
rect 268334 252517 268394 471955
rect 270814 452454 271394 487898
rect 270814 452218 270986 452454
rect 271222 452218 271394 452454
rect 270814 452134 271394 452218
rect 270814 451898 270986 452134
rect 271222 451898 271394 452134
rect 270814 416454 271394 451898
rect 270814 416218 270986 416454
rect 271222 416218 271394 416454
rect 270814 416134 271394 416218
rect 270814 415898 270986 416134
rect 271222 415898 271394 416134
rect 270814 380454 271394 415898
rect 270814 380218 270986 380454
rect 271222 380218 271394 380454
rect 270814 380134 271394 380218
rect 270814 379898 270986 380134
rect 271222 379898 271394 380134
rect 268886 360858 268946 363342
rect 270814 344454 271394 379898
rect 270814 344218 270986 344454
rect 271222 344218 271394 344454
rect 270814 344134 271394 344218
rect 270814 343898 270986 344134
rect 271222 343898 271394 344134
rect 270814 308454 271394 343898
rect 270814 308218 270986 308454
rect 271222 308218 271394 308454
rect 270814 308134 271394 308218
rect 270814 307898 270986 308134
rect 271222 307898 271394 308134
rect 270814 272454 271394 307898
rect 270814 272218 270986 272454
rect 271222 272218 271394 272454
rect 270814 272134 271394 272218
rect 270814 271898 270986 272134
rect 271222 271898 271394 272134
rect 268331 252516 268397 252517
rect 268331 252452 268332 252516
rect 268396 252452 268397 252516
rect 268331 252451 268397 252452
rect 263254 228658 263426 228894
rect 263662 228658 263834 228894
rect 263254 228574 263834 228658
rect 263254 228338 263426 228574
rect 263662 228338 263834 228574
rect 263254 192894 263834 228338
rect 263254 192658 263426 192894
rect 263662 192658 263834 192894
rect 263254 192574 263834 192658
rect 263254 192338 263426 192574
rect 263662 192338 263834 192574
rect 263254 156894 263834 192338
rect 263254 156658 263426 156894
rect 263662 156658 263834 156894
rect 263254 156574 263834 156658
rect 263254 156338 263426 156574
rect 263662 156338 263834 156574
rect 263254 120894 263834 156338
rect 263254 120658 263426 120894
rect 263662 120658 263834 120894
rect 263254 120574 263834 120658
rect 263254 120338 263426 120574
rect 263662 120338 263834 120574
rect 263254 84894 263834 120338
rect 263254 84658 263426 84894
rect 263662 84658 263834 84894
rect 263254 84574 263834 84658
rect 263254 84338 263426 84574
rect 263662 84338 263834 84574
rect 263254 48894 263834 84338
rect 263254 48658 263426 48894
rect 263662 48658 263834 48894
rect 263254 48574 263834 48658
rect 263254 48338 263426 48574
rect 263662 48338 263834 48574
rect 263254 12894 263834 48338
rect 263254 12658 263426 12894
rect 263662 12658 263834 12894
rect 263254 12574 263834 12658
rect 263254 12338 263426 12574
rect 263662 12338 263834 12574
rect 245254 -7022 245426 -6786
rect 245662 -7022 245834 -6786
rect 245254 -7106 245834 -7022
rect 245254 -7342 245426 -7106
rect 245662 -7342 245834 -7106
rect 245254 -7354 245834 -7342
rect 263254 -5866 263834 12338
rect 270814 236454 271394 271898
rect 270814 236218 270986 236454
rect 271222 236218 271394 236454
rect 270814 236134 271394 236218
rect 270814 235898 270986 236134
rect 271222 235898 271394 236134
rect 270814 200454 271394 235898
rect 270814 200218 270986 200454
rect 271222 200218 271394 200454
rect 270814 200134 271394 200218
rect 270814 199898 270986 200134
rect 271222 199898 271394 200134
rect 270814 164454 271394 199898
rect 270814 164218 270986 164454
rect 271222 164218 271394 164454
rect 270814 164134 271394 164218
rect 270814 163898 270986 164134
rect 271222 163898 271394 164134
rect 270814 128454 271394 163898
rect 270814 128218 270986 128454
rect 271222 128218 271394 128454
rect 270814 128134 271394 128218
rect 270814 127898 270986 128134
rect 271222 127898 271394 128134
rect 270814 92454 271394 127898
rect 270814 92218 270986 92454
rect 271222 92218 271394 92454
rect 270814 92134 271394 92218
rect 270814 91898 270986 92134
rect 271222 91898 271394 92134
rect 270814 56454 271394 91898
rect 270814 56218 270986 56454
rect 271222 56218 271394 56454
rect 270814 56134 271394 56218
rect 270814 55898 270986 56134
rect 271222 55898 271394 56134
rect 270814 20454 271394 55898
rect 270814 20218 270986 20454
rect 271222 20218 271394 20454
rect 270814 20134 271394 20218
rect 270814 19898 270986 20134
rect 271222 19898 271394 20134
rect 270814 -1266 271394 19898
rect 270814 -1502 270986 -1266
rect 271222 -1502 271394 -1266
rect 270814 -1586 271394 -1502
rect 270814 -1822 270986 -1586
rect 271222 -1822 271394 -1586
rect 270814 -1834 271394 -1822
rect 274294 671934 274874 707042
rect 274294 671698 274466 671934
rect 274702 671698 274874 671934
rect 274294 671614 274874 671698
rect 274294 671378 274466 671614
rect 274702 671378 274874 671614
rect 274294 635934 274874 671378
rect 274294 635698 274466 635934
rect 274702 635698 274874 635934
rect 274294 635614 274874 635698
rect 274294 635378 274466 635614
rect 274702 635378 274874 635614
rect 274294 599934 274874 635378
rect 274294 599698 274466 599934
rect 274702 599698 274874 599934
rect 274294 599614 274874 599698
rect 274294 599378 274466 599614
rect 274702 599378 274874 599614
rect 274294 563934 274874 599378
rect 274294 563698 274466 563934
rect 274702 563698 274874 563934
rect 274294 563614 274874 563698
rect 274294 563378 274466 563614
rect 274702 563378 274874 563614
rect 274294 527934 274874 563378
rect 274294 527698 274466 527934
rect 274702 527698 274874 527934
rect 274294 527614 274874 527698
rect 274294 527378 274466 527614
rect 274702 527378 274874 527614
rect 274294 491934 274874 527378
rect 274294 491698 274466 491934
rect 274702 491698 274874 491934
rect 274294 491614 274874 491698
rect 274294 491378 274466 491614
rect 274702 491378 274874 491614
rect 274294 455934 274874 491378
rect 274294 455698 274466 455934
rect 274702 455698 274874 455934
rect 274294 455614 274874 455698
rect 274294 455378 274466 455614
rect 274702 455378 274874 455614
rect 274294 419934 274874 455378
rect 274294 419698 274466 419934
rect 274702 419698 274874 419934
rect 274294 419614 274874 419698
rect 274294 419378 274466 419614
rect 274702 419378 274874 419614
rect 274294 383934 274874 419378
rect 274294 383698 274466 383934
rect 274702 383698 274874 383934
rect 274294 383614 274874 383698
rect 274294 383378 274466 383614
rect 274702 383378 274874 383614
rect 274294 347934 274874 383378
rect 274294 347698 274466 347934
rect 274702 347698 274874 347934
rect 274294 347614 274874 347698
rect 274294 347378 274466 347614
rect 274702 347378 274874 347614
rect 274294 311934 274874 347378
rect 274294 311698 274466 311934
rect 274702 311698 274874 311934
rect 274294 311614 274874 311698
rect 274294 311378 274466 311614
rect 274702 311378 274874 311614
rect 274294 275934 274874 311378
rect 274294 275698 274466 275934
rect 274702 275698 274874 275934
rect 274294 275614 274874 275698
rect 274294 275378 274466 275614
rect 274702 275378 274874 275614
rect 274294 239934 274874 275378
rect 274294 239698 274466 239934
rect 274702 239698 274874 239934
rect 274294 239614 274874 239698
rect 274294 239378 274466 239614
rect 274702 239378 274874 239614
rect 274294 203934 274874 239378
rect 274294 203698 274466 203934
rect 274702 203698 274874 203934
rect 274294 203614 274874 203698
rect 274294 203378 274466 203614
rect 274702 203378 274874 203614
rect 274294 167934 274874 203378
rect 274294 167698 274466 167934
rect 274702 167698 274874 167934
rect 274294 167614 274874 167698
rect 274294 167378 274466 167614
rect 274702 167378 274874 167614
rect 274294 131934 274874 167378
rect 274294 131698 274466 131934
rect 274702 131698 274874 131934
rect 274294 131614 274874 131698
rect 274294 131378 274466 131614
rect 274702 131378 274874 131614
rect 274294 95934 274874 131378
rect 274294 95698 274466 95934
rect 274702 95698 274874 95934
rect 274294 95614 274874 95698
rect 274294 95378 274466 95614
rect 274702 95378 274874 95614
rect 274294 59934 274874 95378
rect 274294 59698 274466 59934
rect 274702 59698 274874 59934
rect 274294 59614 274874 59698
rect 274294 59378 274466 59614
rect 274702 59378 274874 59614
rect 274294 23934 274874 59378
rect 274294 23698 274466 23934
rect 274702 23698 274874 23934
rect 274294 23614 274874 23698
rect 274294 23378 274466 23614
rect 274702 23378 274874 23614
rect 274294 -3106 274874 23378
rect 274294 -3342 274466 -3106
rect 274702 -3342 274874 -3106
rect 274294 -3426 274874 -3342
rect 274294 -3662 274466 -3426
rect 274702 -3662 274874 -3426
rect 274294 -3674 274874 -3662
rect 277774 675414 278354 708882
rect 277774 675178 277946 675414
rect 278182 675178 278354 675414
rect 277774 675094 278354 675178
rect 277774 674858 277946 675094
rect 278182 674858 278354 675094
rect 277774 639414 278354 674858
rect 277774 639178 277946 639414
rect 278182 639178 278354 639414
rect 277774 639094 278354 639178
rect 277774 638858 277946 639094
rect 278182 638858 278354 639094
rect 277774 603414 278354 638858
rect 277774 603178 277946 603414
rect 278182 603178 278354 603414
rect 277774 603094 278354 603178
rect 277774 602858 277946 603094
rect 278182 602858 278354 603094
rect 277774 567414 278354 602858
rect 277774 567178 277946 567414
rect 278182 567178 278354 567414
rect 277774 567094 278354 567178
rect 277774 566858 277946 567094
rect 278182 566858 278354 567094
rect 277774 531414 278354 566858
rect 277774 531178 277946 531414
rect 278182 531178 278354 531414
rect 277774 531094 278354 531178
rect 277774 530858 277946 531094
rect 278182 530858 278354 531094
rect 277774 495414 278354 530858
rect 277774 495178 277946 495414
rect 278182 495178 278354 495414
rect 277774 495094 278354 495178
rect 277774 494858 277946 495094
rect 278182 494858 278354 495094
rect 277774 459414 278354 494858
rect 277774 459178 277946 459414
rect 278182 459178 278354 459414
rect 277774 459094 278354 459178
rect 277774 458858 277946 459094
rect 278182 458858 278354 459094
rect 277774 423414 278354 458858
rect 277774 423178 277946 423414
rect 278182 423178 278354 423414
rect 277774 423094 278354 423178
rect 277774 422858 277946 423094
rect 278182 422858 278354 423094
rect 277774 387414 278354 422858
rect 277774 387178 277946 387414
rect 278182 387178 278354 387414
rect 277774 387094 278354 387178
rect 277774 386858 277946 387094
rect 278182 386858 278354 387094
rect 277774 351414 278354 386858
rect 277774 351178 277946 351414
rect 278182 351178 278354 351414
rect 277774 351094 278354 351178
rect 277774 350858 277946 351094
rect 278182 350858 278354 351094
rect 277774 315414 278354 350858
rect 277774 315178 277946 315414
rect 278182 315178 278354 315414
rect 277774 315094 278354 315178
rect 277774 314858 277946 315094
rect 278182 314858 278354 315094
rect 277774 279414 278354 314858
rect 277774 279178 277946 279414
rect 278182 279178 278354 279414
rect 277774 279094 278354 279178
rect 277774 278858 277946 279094
rect 278182 278858 278354 279094
rect 277774 243414 278354 278858
rect 277774 243178 277946 243414
rect 278182 243178 278354 243414
rect 277774 243094 278354 243178
rect 277774 242858 277946 243094
rect 278182 242858 278354 243094
rect 277774 207414 278354 242858
rect 277774 207178 277946 207414
rect 278182 207178 278354 207414
rect 277774 207094 278354 207178
rect 277774 206858 277946 207094
rect 278182 206858 278354 207094
rect 277774 171414 278354 206858
rect 277774 171178 277946 171414
rect 278182 171178 278354 171414
rect 277774 171094 278354 171178
rect 277774 170858 277946 171094
rect 278182 170858 278354 171094
rect 277774 135414 278354 170858
rect 277774 135178 277946 135414
rect 278182 135178 278354 135414
rect 277774 135094 278354 135178
rect 277774 134858 277946 135094
rect 278182 134858 278354 135094
rect 277774 99414 278354 134858
rect 277774 99178 277946 99414
rect 278182 99178 278354 99414
rect 277774 99094 278354 99178
rect 277774 98858 277946 99094
rect 278182 98858 278354 99094
rect 277774 63414 278354 98858
rect 277774 63178 277946 63414
rect 278182 63178 278354 63414
rect 277774 63094 278354 63178
rect 277774 62858 277946 63094
rect 278182 62858 278354 63094
rect 277774 27414 278354 62858
rect 277774 27178 277946 27414
rect 278182 27178 278354 27414
rect 277774 27094 278354 27178
rect 277774 26858 277946 27094
rect 278182 26858 278354 27094
rect 277774 -4946 278354 26858
rect 277774 -5182 277946 -4946
rect 278182 -5182 278354 -4946
rect 277774 -5266 278354 -5182
rect 277774 -5502 277946 -5266
rect 278182 -5502 278354 -5266
rect 277774 -5514 278354 -5502
rect 281254 678894 281834 710722
rect 299254 710358 299834 711290
rect 299254 710122 299426 710358
rect 299662 710122 299834 710358
rect 299254 710038 299834 710122
rect 299254 709802 299426 710038
rect 299662 709802 299834 710038
rect 295774 708518 296354 709450
rect 295774 708282 295946 708518
rect 296182 708282 296354 708518
rect 295774 708198 296354 708282
rect 295774 707962 295946 708198
rect 296182 707962 296354 708198
rect 292294 706678 292874 707610
rect 292294 706442 292466 706678
rect 292702 706442 292874 706678
rect 292294 706358 292874 706442
rect 292294 706122 292466 706358
rect 292702 706122 292874 706358
rect 281254 678658 281426 678894
rect 281662 678658 281834 678894
rect 281254 678574 281834 678658
rect 281254 678338 281426 678574
rect 281662 678338 281834 678574
rect 281254 642894 281834 678338
rect 281254 642658 281426 642894
rect 281662 642658 281834 642894
rect 281254 642574 281834 642658
rect 281254 642338 281426 642574
rect 281662 642338 281834 642574
rect 281254 606894 281834 642338
rect 281254 606658 281426 606894
rect 281662 606658 281834 606894
rect 281254 606574 281834 606658
rect 281254 606338 281426 606574
rect 281662 606338 281834 606574
rect 281254 570894 281834 606338
rect 281254 570658 281426 570894
rect 281662 570658 281834 570894
rect 281254 570574 281834 570658
rect 281254 570338 281426 570574
rect 281662 570338 281834 570574
rect 281254 534894 281834 570338
rect 281254 534658 281426 534894
rect 281662 534658 281834 534894
rect 281254 534574 281834 534658
rect 281254 534338 281426 534574
rect 281662 534338 281834 534574
rect 281254 498894 281834 534338
rect 281254 498658 281426 498894
rect 281662 498658 281834 498894
rect 281254 498574 281834 498658
rect 281254 498338 281426 498574
rect 281662 498338 281834 498574
rect 281254 462894 281834 498338
rect 281254 462658 281426 462894
rect 281662 462658 281834 462894
rect 281254 462574 281834 462658
rect 281254 462338 281426 462574
rect 281662 462338 281834 462574
rect 281254 426894 281834 462338
rect 281254 426658 281426 426894
rect 281662 426658 281834 426894
rect 281254 426574 281834 426658
rect 281254 426338 281426 426574
rect 281662 426338 281834 426574
rect 281254 390894 281834 426338
rect 281254 390658 281426 390894
rect 281662 390658 281834 390894
rect 281254 390574 281834 390658
rect 281254 390338 281426 390574
rect 281662 390338 281834 390574
rect 281254 354894 281834 390338
rect 281254 354658 281426 354894
rect 281662 354658 281834 354894
rect 281254 354574 281834 354658
rect 281254 354338 281426 354574
rect 281662 354338 281834 354574
rect 281254 318894 281834 354338
rect 281254 318658 281426 318894
rect 281662 318658 281834 318894
rect 281254 318574 281834 318658
rect 281254 318338 281426 318574
rect 281662 318338 281834 318574
rect 281254 282894 281834 318338
rect 281254 282658 281426 282894
rect 281662 282658 281834 282894
rect 281254 282574 281834 282658
rect 281254 282338 281426 282574
rect 281662 282338 281834 282574
rect 281254 246894 281834 282338
rect 281254 246658 281426 246894
rect 281662 246658 281834 246894
rect 281254 246574 281834 246658
rect 281254 246338 281426 246574
rect 281662 246338 281834 246574
rect 281254 210894 281834 246338
rect 281254 210658 281426 210894
rect 281662 210658 281834 210894
rect 281254 210574 281834 210658
rect 281254 210338 281426 210574
rect 281662 210338 281834 210574
rect 281254 174894 281834 210338
rect 281254 174658 281426 174894
rect 281662 174658 281834 174894
rect 281254 174574 281834 174658
rect 281254 174338 281426 174574
rect 281662 174338 281834 174574
rect 281254 138894 281834 174338
rect 281254 138658 281426 138894
rect 281662 138658 281834 138894
rect 281254 138574 281834 138658
rect 281254 138338 281426 138574
rect 281662 138338 281834 138574
rect 281254 102894 281834 138338
rect 281254 102658 281426 102894
rect 281662 102658 281834 102894
rect 281254 102574 281834 102658
rect 281254 102338 281426 102574
rect 281662 102338 281834 102574
rect 281254 66894 281834 102338
rect 281254 66658 281426 66894
rect 281662 66658 281834 66894
rect 281254 66574 281834 66658
rect 281254 66338 281426 66574
rect 281662 66338 281834 66574
rect 281254 30894 281834 66338
rect 281254 30658 281426 30894
rect 281662 30658 281834 30894
rect 281254 30574 281834 30658
rect 281254 30338 281426 30574
rect 281662 30338 281834 30574
rect 263254 -6102 263426 -5866
rect 263662 -6102 263834 -5866
rect 263254 -6186 263834 -6102
rect 263254 -6422 263426 -6186
rect 263662 -6422 263834 -6186
rect 263254 -7354 263834 -6422
rect 281254 -6786 281834 30338
rect 288814 704838 289394 705770
rect 288814 704602 288986 704838
rect 289222 704602 289394 704838
rect 288814 704518 289394 704602
rect 288814 704282 288986 704518
rect 289222 704282 289394 704518
rect 288814 686454 289394 704282
rect 288814 686218 288986 686454
rect 289222 686218 289394 686454
rect 288814 686134 289394 686218
rect 288814 685898 288986 686134
rect 289222 685898 289394 686134
rect 288814 650454 289394 685898
rect 288814 650218 288986 650454
rect 289222 650218 289394 650454
rect 288814 650134 289394 650218
rect 288814 649898 288986 650134
rect 289222 649898 289394 650134
rect 288814 614454 289394 649898
rect 288814 614218 288986 614454
rect 289222 614218 289394 614454
rect 288814 614134 289394 614218
rect 288814 613898 288986 614134
rect 289222 613898 289394 614134
rect 288814 578454 289394 613898
rect 288814 578218 288986 578454
rect 289222 578218 289394 578454
rect 288814 578134 289394 578218
rect 288814 577898 288986 578134
rect 289222 577898 289394 578134
rect 288814 542454 289394 577898
rect 288814 542218 288986 542454
rect 289222 542218 289394 542454
rect 288814 542134 289394 542218
rect 288814 541898 288986 542134
rect 289222 541898 289394 542134
rect 288814 506454 289394 541898
rect 288814 506218 288986 506454
rect 289222 506218 289394 506454
rect 288814 506134 289394 506218
rect 288814 505898 288986 506134
rect 289222 505898 289394 506134
rect 288814 470454 289394 505898
rect 288814 470218 288986 470454
rect 289222 470218 289394 470454
rect 288814 470134 289394 470218
rect 288814 469898 288986 470134
rect 289222 469898 289394 470134
rect 288814 434454 289394 469898
rect 288814 434218 288986 434454
rect 289222 434218 289394 434454
rect 288814 434134 289394 434218
rect 288814 433898 288986 434134
rect 289222 433898 289394 434134
rect 288814 398454 289394 433898
rect 288814 398218 288986 398454
rect 289222 398218 289394 398454
rect 288814 398134 289394 398218
rect 288814 397898 288986 398134
rect 289222 397898 289394 398134
rect 288814 362454 289394 397898
rect 288814 362218 288986 362454
rect 289222 362218 289394 362454
rect 288814 362134 289394 362218
rect 288814 361898 288986 362134
rect 289222 361898 289394 362134
rect 288814 326454 289394 361898
rect 288814 326218 288986 326454
rect 289222 326218 289394 326454
rect 288814 326134 289394 326218
rect 288814 325898 288986 326134
rect 289222 325898 289394 326134
rect 288814 290454 289394 325898
rect 288814 290218 288986 290454
rect 289222 290218 289394 290454
rect 288814 290134 289394 290218
rect 288814 289898 288986 290134
rect 289222 289898 289394 290134
rect 288814 254454 289394 289898
rect 288814 254218 288986 254454
rect 289222 254218 289394 254454
rect 288814 254134 289394 254218
rect 288814 253898 288986 254134
rect 289222 253898 289394 254134
rect 288814 218454 289394 253898
rect 288814 218218 288986 218454
rect 289222 218218 289394 218454
rect 288814 218134 289394 218218
rect 288814 217898 288986 218134
rect 289222 217898 289394 218134
rect 288814 182454 289394 217898
rect 288814 182218 288986 182454
rect 289222 182218 289394 182454
rect 288814 182134 289394 182218
rect 288814 181898 288986 182134
rect 289222 181898 289394 182134
rect 288814 146454 289394 181898
rect 288814 146218 288986 146454
rect 289222 146218 289394 146454
rect 288814 146134 289394 146218
rect 288814 145898 288986 146134
rect 289222 145898 289394 146134
rect 288814 110454 289394 145898
rect 288814 110218 288986 110454
rect 289222 110218 289394 110454
rect 288814 110134 289394 110218
rect 288814 109898 288986 110134
rect 289222 109898 289394 110134
rect 288814 74454 289394 109898
rect 288814 74218 288986 74454
rect 289222 74218 289394 74454
rect 288814 74134 289394 74218
rect 288814 73898 288986 74134
rect 289222 73898 289394 74134
rect 288814 38454 289394 73898
rect 288814 38218 288986 38454
rect 289222 38218 289394 38454
rect 288814 38134 289394 38218
rect 288814 37898 288986 38134
rect 289222 37898 289394 38134
rect 288814 2454 289394 37898
rect 288814 2218 288986 2454
rect 289222 2218 289394 2454
rect 288814 2134 289394 2218
rect 288814 1898 288986 2134
rect 289222 1898 289394 2134
rect 288814 -346 289394 1898
rect 288814 -582 288986 -346
rect 289222 -582 289394 -346
rect 288814 -666 289394 -582
rect 288814 -902 288986 -666
rect 289222 -902 289394 -666
rect 288814 -1834 289394 -902
rect 292294 689934 292874 706122
rect 292294 689698 292466 689934
rect 292702 689698 292874 689934
rect 292294 689614 292874 689698
rect 292294 689378 292466 689614
rect 292702 689378 292874 689614
rect 292294 653934 292874 689378
rect 292294 653698 292466 653934
rect 292702 653698 292874 653934
rect 292294 653614 292874 653698
rect 292294 653378 292466 653614
rect 292702 653378 292874 653614
rect 292294 617934 292874 653378
rect 292294 617698 292466 617934
rect 292702 617698 292874 617934
rect 292294 617614 292874 617698
rect 292294 617378 292466 617614
rect 292702 617378 292874 617614
rect 292294 581934 292874 617378
rect 292294 581698 292466 581934
rect 292702 581698 292874 581934
rect 292294 581614 292874 581698
rect 292294 581378 292466 581614
rect 292702 581378 292874 581614
rect 292294 545934 292874 581378
rect 292294 545698 292466 545934
rect 292702 545698 292874 545934
rect 292294 545614 292874 545698
rect 292294 545378 292466 545614
rect 292702 545378 292874 545614
rect 292294 509934 292874 545378
rect 292294 509698 292466 509934
rect 292702 509698 292874 509934
rect 292294 509614 292874 509698
rect 292294 509378 292466 509614
rect 292702 509378 292874 509614
rect 292294 473934 292874 509378
rect 292294 473698 292466 473934
rect 292702 473698 292874 473934
rect 292294 473614 292874 473698
rect 292294 473378 292466 473614
rect 292702 473378 292874 473614
rect 292294 437934 292874 473378
rect 292294 437698 292466 437934
rect 292702 437698 292874 437934
rect 292294 437614 292874 437698
rect 292294 437378 292466 437614
rect 292702 437378 292874 437614
rect 292294 401934 292874 437378
rect 292294 401698 292466 401934
rect 292702 401698 292874 401934
rect 292294 401614 292874 401698
rect 292294 401378 292466 401614
rect 292702 401378 292874 401614
rect 292294 365934 292874 401378
rect 292294 365698 292466 365934
rect 292702 365698 292874 365934
rect 292294 365614 292874 365698
rect 292294 365378 292466 365614
rect 292702 365378 292874 365614
rect 292294 329934 292874 365378
rect 292294 329698 292466 329934
rect 292702 329698 292874 329934
rect 292294 329614 292874 329698
rect 292294 329378 292466 329614
rect 292702 329378 292874 329614
rect 292294 293934 292874 329378
rect 292294 293698 292466 293934
rect 292702 293698 292874 293934
rect 292294 293614 292874 293698
rect 292294 293378 292466 293614
rect 292702 293378 292874 293614
rect 292294 257934 292874 293378
rect 292294 257698 292466 257934
rect 292702 257698 292874 257934
rect 292294 257614 292874 257698
rect 292294 257378 292466 257614
rect 292702 257378 292874 257614
rect 292294 221934 292874 257378
rect 292294 221698 292466 221934
rect 292702 221698 292874 221934
rect 292294 221614 292874 221698
rect 292294 221378 292466 221614
rect 292702 221378 292874 221614
rect 292294 185934 292874 221378
rect 292294 185698 292466 185934
rect 292702 185698 292874 185934
rect 292294 185614 292874 185698
rect 292294 185378 292466 185614
rect 292702 185378 292874 185614
rect 292294 149934 292874 185378
rect 292294 149698 292466 149934
rect 292702 149698 292874 149934
rect 292294 149614 292874 149698
rect 292294 149378 292466 149614
rect 292702 149378 292874 149614
rect 292294 113934 292874 149378
rect 292294 113698 292466 113934
rect 292702 113698 292874 113934
rect 292294 113614 292874 113698
rect 292294 113378 292466 113614
rect 292702 113378 292874 113614
rect 292294 77934 292874 113378
rect 292294 77698 292466 77934
rect 292702 77698 292874 77934
rect 292294 77614 292874 77698
rect 292294 77378 292466 77614
rect 292702 77378 292874 77614
rect 292294 41934 292874 77378
rect 292294 41698 292466 41934
rect 292702 41698 292874 41934
rect 292294 41614 292874 41698
rect 292294 41378 292466 41614
rect 292702 41378 292874 41614
rect 292294 5934 292874 41378
rect 292294 5698 292466 5934
rect 292702 5698 292874 5934
rect 292294 5614 292874 5698
rect 292294 5378 292466 5614
rect 292702 5378 292874 5614
rect 292294 -2186 292874 5378
rect 292294 -2422 292466 -2186
rect 292702 -2422 292874 -2186
rect 292294 -2506 292874 -2422
rect 292294 -2742 292466 -2506
rect 292702 -2742 292874 -2506
rect 292294 -3674 292874 -2742
rect 295774 693414 296354 707962
rect 295774 693178 295946 693414
rect 296182 693178 296354 693414
rect 295774 693094 296354 693178
rect 295774 692858 295946 693094
rect 296182 692858 296354 693094
rect 295774 657414 296354 692858
rect 295774 657178 295946 657414
rect 296182 657178 296354 657414
rect 295774 657094 296354 657178
rect 295774 656858 295946 657094
rect 296182 656858 296354 657094
rect 295774 621414 296354 656858
rect 295774 621178 295946 621414
rect 296182 621178 296354 621414
rect 295774 621094 296354 621178
rect 295774 620858 295946 621094
rect 296182 620858 296354 621094
rect 295774 585414 296354 620858
rect 295774 585178 295946 585414
rect 296182 585178 296354 585414
rect 295774 585094 296354 585178
rect 295774 584858 295946 585094
rect 296182 584858 296354 585094
rect 295774 549414 296354 584858
rect 295774 549178 295946 549414
rect 296182 549178 296354 549414
rect 295774 549094 296354 549178
rect 295774 548858 295946 549094
rect 296182 548858 296354 549094
rect 295774 513414 296354 548858
rect 295774 513178 295946 513414
rect 296182 513178 296354 513414
rect 295774 513094 296354 513178
rect 295774 512858 295946 513094
rect 296182 512858 296354 513094
rect 295774 477414 296354 512858
rect 295774 477178 295946 477414
rect 296182 477178 296354 477414
rect 295774 477094 296354 477178
rect 295774 476858 295946 477094
rect 296182 476858 296354 477094
rect 295774 441414 296354 476858
rect 295774 441178 295946 441414
rect 296182 441178 296354 441414
rect 295774 441094 296354 441178
rect 295774 440858 295946 441094
rect 296182 440858 296354 441094
rect 295774 405414 296354 440858
rect 295774 405178 295946 405414
rect 296182 405178 296354 405414
rect 295774 405094 296354 405178
rect 295774 404858 295946 405094
rect 296182 404858 296354 405094
rect 295774 369414 296354 404858
rect 295774 369178 295946 369414
rect 296182 369178 296354 369414
rect 295774 369094 296354 369178
rect 295774 368858 295946 369094
rect 296182 368858 296354 369094
rect 295774 333414 296354 368858
rect 295774 333178 295946 333414
rect 296182 333178 296354 333414
rect 295774 333094 296354 333178
rect 295774 332858 295946 333094
rect 296182 332858 296354 333094
rect 295774 297414 296354 332858
rect 295774 297178 295946 297414
rect 296182 297178 296354 297414
rect 295774 297094 296354 297178
rect 295774 296858 295946 297094
rect 296182 296858 296354 297094
rect 295774 261414 296354 296858
rect 295774 261178 295946 261414
rect 296182 261178 296354 261414
rect 295774 261094 296354 261178
rect 295774 260858 295946 261094
rect 296182 260858 296354 261094
rect 295774 225414 296354 260858
rect 295774 225178 295946 225414
rect 296182 225178 296354 225414
rect 295774 225094 296354 225178
rect 295774 224858 295946 225094
rect 296182 224858 296354 225094
rect 295774 189414 296354 224858
rect 295774 189178 295946 189414
rect 296182 189178 296354 189414
rect 295774 189094 296354 189178
rect 295774 188858 295946 189094
rect 296182 188858 296354 189094
rect 295774 153414 296354 188858
rect 295774 153178 295946 153414
rect 296182 153178 296354 153414
rect 295774 153094 296354 153178
rect 295774 152858 295946 153094
rect 296182 152858 296354 153094
rect 295774 117414 296354 152858
rect 295774 117178 295946 117414
rect 296182 117178 296354 117414
rect 295774 117094 296354 117178
rect 295774 116858 295946 117094
rect 296182 116858 296354 117094
rect 295774 81414 296354 116858
rect 295774 81178 295946 81414
rect 296182 81178 296354 81414
rect 295774 81094 296354 81178
rect 295774 80858 295946 81094
rect 296182 80858 296354 81094
rect 295774 45414 296354 80858
rect 295774 45178 295946 45414
rect 296182 45178 296354 45414
rect 295774 45094 296354 45178
rect 295774 44858 295946 45094
rect 296182 44858 296354 45094
rect 295774 9414 296354 44858
rect 295774 9178 295946 9414
rect 296182 9178 296354 9414
rect 295774 9094 296354 9178
rect 295774 8858 295946 9094
rect 296182 8858 296354 9094
rect 295774 -4026 296354 8858
rect 295774 -4262 295946 -4026
rect 296182 -4262 296354 -4026
rect 295774 -4346 296354 -4262
rect 295774 -4582 295946 -4346
rect 296182 -4582 296354 -4346
rect 295774 -5514 296354 -4582
rect 299254 696894 299834 709802
rect 317254 711278 317834 711290
rect 317254 711042 317426 711278
rect 317662 711042 317834 711278
rect 317254 710958 317834 711042
rect 317254 710722 317426 710958
rect 317662 710722 317834 710958
rect 313774 709438 314354 709450
rect 313774 709202 313946 709438
rect 314182 709202 314354 709438
rect 313774 709118 314354 709202
rect 313774 708882 313946 709118
rect 314182 708882 314354 709118
rect 310294 707598 310874 707610
rect 310294 707362 310466 707598
rect 310702 707362 310874 707598
rect 310294 707278 310874 707362
rect 310294 707042 310466 707278
rect 310702 707042 310874 707278
rect 299254 696658 299426 696894
rect 299662 696658 299834 696894
rect 299254 696574 299834 696658
rect 299254 696338 299426 696574
rect 299662 696338 299834 696574
rect 299254 660894 299834 696338
rect 299254 660658 299426 660894
rect 299662 660658 299834 660894
rect 299254 660574 299834 660658
rect 299254 660338 299426 660574
rect 299662 660338 299834 660574
rect 299254 624894 299834 660338
rect 299254 624658 299426 624894
rect 299662 624658 299834 624894
rect 299254 624574 299834 624658
rect 299254 624338 299426 624574
rect 299662 624338 299834 624574
rect 299254 588894 299834 624338
rect 299254 588658 299426 588894
rect 299662 588658 299834 588894
rect 299254 588574 299834 588658
rect 299254 588338 299426 588574
rect 299662 588338 299834 588574
rect 299254 552894 299834 588338
rect 299254 552658 299426 552894
rect 299662 552658 299834 552894
rect 299254 552574 299834 552658
rect 299254 552338 299426 552574
rect 299662 552338 299834 552574
rect 299254 516894 299834 552338
rect 299254 516658 299426 516894
rect 299662 516658 299834 516894
rect 299254 516574 299834 516658
rect 299254 516338 299426 516574
rect 299662 516338 299834 516574
rect 299254 480894 299834 516338
rect 299254 480658 299426 480894
rect 299662 480658 299834 480894
rect 299254 480574 299834 480658
rect 299254 480338 299426 480574
rect 299662 480338 299834 480574
rect 299254 444894 299834 480338
rect 299254 444658 299426 444894
rect 299662 444658 299834 444894
rect 299254 444574 299834 444658
rect 299254 444338 299426 444574
rect 299662 444338 299834 444574
rect 299254 408894 299834 444338
rect 299254 408658 299426 408894
rect 299662 408658 299834 408894
rect 299254 408574 299834 408658
rect 299254 408338 299426 408574
rect 299662 408338 299834 408574
rect 299254 372894 299834 408338
rect 299254 372658 299426 372894
rect 299662 372658 299834 372894
rect 299254 372574 299834 372658
rect 299254 372338 299426 372574
rect 299662 372338 299834 372574
rect 299254 336894 299834 372338
rect 299254 336658 299426 336894
rect 299662 336658 299834 336894
rect 299254 336574 299834 336658
rect 299254 336338 299426 336574
rect 299662 336338 299834 336574
rect 299254 300894 299834 336338
rect 299254 300658 299426 300894
rect 299662 300658 299834 300894
rect 299254 300574 299834 300658
rect 299254 300338 299426 300574
rect 299662 300338 299834 300574
rect 299254 264894 299834 300338
rect 299254 264658 299426 264894
rect 299662 264658 299834 264894
rect 299254 264574 299834 264658
rect 299254 264338 299426 264574
rect 299662 264338 299834 264574
rect 299254 228894 299834 264338
rect 299254 228658 299426 228894
rect 299662 228658 299834 228894
rect 299254 228574 299834 228658
rect 299254 228338 299426 228574
rect 299662 228338 299834 228574
rect 299254 192894 299834 228338
rect 299254 192658 299426 192894
rect 299662 192658 299834 192894
rect 299254 192574 299834 192658
rect 299254 192338 299426 192574
rect 299662 192338 299834 192574
rect 299254 156894 299834 192338
rect 299254 156658 299426 156894
rect 299662 156658 299834 156894
rect 299254 156574 299834 156658
rect 299254 156338 299426 156574
rect 299662 156338 299834 156574
rect 299254 120894 299834 156338
rect 299254 120658 299426 120894
rect 299662 120658 299834 120894
rect 299254 120574 299834 120658
rect 299254 120338 299426 120574
rect 299662 120338 299834 120574
rect 299254 84894 299834 120338
rect 299254 84658 299426 84894
rect 299662 84658 299834 84894
rect 299254 84574 299834 84658
rect 299254 84338 299426 84574
rect 299662 84338 299834 84574
rect 299254 48894 299834 84338
rect 299254 48658 299426 48894
rect 299662 48658 299834 48894
rect 299254 48574 299834 48658
rect 299254 48338 299426 48574
rect 299662 48338 299834 48574
rect 299254 12894 299834 48338
rect 299254 12658 299426 12894
rect 299662 12658 299834 12894
rect 299254 12574 299834 12658
rect 299254 12338 299426 12574
rect 299662 12338 299834 12574
rect 281254 -7022 281426 -6786
rect 281662 -7022 281834 -6786
rect 281254 -7106 281834 -7022
rect 281254 -7342 281426 -7106
rect 281662 -7342 281834 -7106
rect 281254 -7354 281834 -7342
rect 299254 -5866 299834 12338
rect 306814 705758 307394 705770
rect 306814 705522 306986 705758
rect 307222 705522 307394 705758
rect 306814 705438 307394 705522
rect 306814 705202 306986 705438
rect 307222 705202 307394 705438
rect 306814 668454 307394 705202
rect 306814 668218 306986 668454
rect 307222 668218 307394 668454
rect 306814 668134 307394 668218
rect 306814 667898 306986 668134
rect 307222 667898 307394 668134
rect 306814 632454 307394 667898
rect 306814 632218 306986 632454
rect 307222 632218 307394 632454
rect 306814 632134 307394 632218
rect 306814 631898 306986 632134
rect 307222 631898 307394 632134
rect 306814 596454 307394 631898
rect 306814 596218 306986 596454
rect 307222 596218 307394 596454
rect 306814 596134 307394 596218
rect 306814 595898 306986 596134
rect 307222 595898 307394 596134
rect 306814 560454 307394 595898
rect 306814 560218 306986 560454
rect 307222 560218 307394 560454
rect 306814 560134 307394 560218
rect 306814 559898 306986 560134
rect 307222 559898 307394 560134
rect 306814 524454 307394 559898
rect 306814 524218 306986 524454
rect 307222 524218 307394 524454
rect 306814 524134 307394 524218
rect 306814 523898 306986 524134
rect 307222 523898 307394 524134
rect 306814 488454 307394 523898
rect 306814 488218 306986 488454
rect 307222 488218 307394 488454
rect 306814 488134 307394 488218
rect 306814 487898 306986 488134
rect 307222 487898 307394 488134
rect 306814 452454 307394 487898
rect 306814 452218 306986 452454
rect 307222 452218 307394 452454
rect 306814 452134 307394 452218
rect 306814 451898 306986 452134
rect 307222 451898 307394 452134
rect 306814 416454 307394 451898
rect 306814 416218 306986 416454
rect 307222 416218 307394 416454
rect 306814 416134 307394 416218
rect 306814 415898 306986 416134
rect 307222 415898 307394 416134
rect 306814 380454 307394 415898
rect 306814 380218 306986 380454
rect 307222 380218 307394 380454
rect 306814 380134 307394 380218
rect 306814 379898 306986 380134
rect 307222 379898 307394 380134
rect 306814 344454 307394 379898
rect 306814 344218 306986 344454
rect 307222 344218 307394 344454
rect 306814 344134 307394 344218
rect 306814 343898 306986 344134
rect 307222 343898 307394 344134
rect 306814 308454 307394 343898
rect 306814 308218 306986 308454
rect 307222 308218 307394 308454
rect 306814 308134 307394 308218
rect 306814 307898 306986 308134
rect 307222 307898 307394 308134
rect 306814 272454 307394 307898
rect 306814 272218 306986 272454
rect 307222 272218 307394 272454
rect 306814 272134 307394 272218
rect 306814 271898 306986 272134
rect 307222 271898 307394 272134
rect 306814 236454 307394 271898
rect 306814 236218 306986 236454
rect 307222 236218 307394 236454
rect 306814 236134 307394 236218
rect 306814 235898 306986 236134
rect 307222 235898 307394 236134
rect 306814 200454 307394 235898
rect 306814 200218 306986 200454
rect 307222 200218 307394 200454
rect 306814 200134 307394 200218
rect 306814 199898 306986 200134
rect 307222 199898 307394 200134
rect 306814 164454 307394 199898
rect 306814 164218 306986 164454
rect 307222 164218 307394 164454
rect 306814 164134 307394 164218
rect 306814 163898 306986 164134
rect 307222 163898 307394 164134
rect 306814 128454 307394 163898
rect 306814 128218 306986 128454
rect 307222 128218 307394 128454
rect 306814 128134 307394 128218
rect 306814 127898 306986 128134
rect 307222 127898 307394 128134
rect 306814 92454 307394 127898
rect 306814 92218 306986 92454
rect 307222 92218 307394 92454
rect 306814 92134 307394 92218
rect 306814 91898 306986 92134
rect 307222 91898 307394 92134
rect 306814 56454 307394 91898
rect 306814 56218 306986 56454
rect 307222 56218 307394 56454
rect 306814 56134 307394 56218
rect 306814 55898 306986 56134
rect 307222 55898 307394 56134
rect 306814 20454 307394 55898
rect 306814 20218 306986 20454
rect 307222 20218 307394 20454
rect 306814 20134 307394 20218
rect 306814 19898 306986 20134
rect 307222 19898 307394 20134
rect 306814 -1266 307394 19898
rect 306814 -1502 306986 -1266
rect 307222 -1502 307394 -1266
rect 306814 -1586 307394 -1502
rect 306814 -1822 306986 -1586
rect 307222 -1822 307394 -1586
rect 306814 -1834 307394 -1822
rect 310294 671934 310874 707042
rect 310294 671698 310466 671934
rect 310702 671698 310874 671934
rect 310294 671614 310874 671698
rect 310294 671378 310466 671614
rect 310702 671378 310874 671614
rect 310294 635934 310874 671378
rect 310294 635698 310466 635934
rect 310702 635698 310874 635934
rect 310294 635614 310874 635698
rect 310294 635378 310466 635614
rect 310702 635378 310874 635614
rect 310294 599934 310874 635378
rect 310294 599698 310466 599934
rect 310702 599698 310874 599934
rect 310294 599614 310874 599698
rect 310294 599378 310466 599614
rect 310702 599378 310874 599614
rect 310294 563934 310874 599378
rect 310294 563698 310466 563934
rect 310702 563698 310874 563934
rect 310294 563614 310874 563698
rect 310294 563378 310466 563614
rect 310702 563378 310874 563614
rect 310294 527934 310874 563378
rect 310294 527698 310466 527934
rect 310702 527698 310874 527934
rect 310294 527614 310874 527698
rect 310294 527378 310466 527614
rect 310702 527378 310874 527614
rect 310294 491934 310874 527378
rect 310294 491698 310466 491934
rect 310702 491698 310874 491934
rect 310294 491614 310874 491698
rect 310294 491378 310466 491614
rect 310702 491378 310874 491614
rect 310294 455934 310874 491378
rect 310294 455698 310466 455934
rect 310702 455698 310874 455934
rect 310294 455614 310874 455698
rect 310294 455378 310466 455614
rect 310702 455378 310874 455614
rect 310294 419934 310874 455378
rect 310294 419698 310466 419934
rect 310702 419698 310874 419934
rect 310294 419614 310874 419698
rect 310294 419378 310466 419614
rect 310702 419378 310874 419614
rect 310294 383934 310874 419378
rect 310294 383698 310466 383934
rect 310702 383698 310874 383934
rect 310294 383614 310874 383698
rect 310294 383378 310466 383614
rect 310702 383378 310874 383614
rect 310294 347934 310874 383378
rect 310294 347698 310466 347934
rect 310702 347698 310874 347934
rect 310294 347614 310874 347698
rect 310294 347378 310466 347614
rect 310702 347378 310874 347614
rect 310294 311934 310874 347378
rect 310294 311698 310466 311934
rect 310702 311698 310874 311934
rect 310294 311614 310874 311698
rect 310294 311378 310466 311614
rect 310702 311378 310874 311614
rect 310294 275934 310874 311378
rect 310294 275698 310466 275934
rect 310702 275698 310874 275934
rect 310294 275614 310874 275698
rect 310294 275378 310466 275614
rect 310702 275378 310874 275614
rect 310294 239934 310874 275378
rect 310294 239698 310466 239934
rect 310702 239698 310874 239934
rect 310294 239614 310874 239698
rect 310294 239378 310466 239614
rect 310702 239378 310874 239614
rect 310294 203934 310874 239378
rect 310294 203698 310466 203934
rect 310702 203698 310874 203934
rect 310294 203614 310874 203698
rect 310294 203378 310466 203614
rect 310702 203378 310874 203614
rect 310294 167934 310874 203378
rect 310294 167698 310466 167934
rect 310702 167698 310874 167934
rect 310294 167614 310874 167698
rect 310294 167378 310466 167614
rect 310702 167378 310874 167614
rect 310294 131934 310874 167378
rect 310294 131698 310466 131934
rect 310702 131698 310874 131934
rect 310294 131614 310874 131698
rect 310294 131378 310466 131614
rect 310702 131378 310874 131614
rect 310294 95934 310874 131378
rect 310294 95698 310466 95934
rect 310702 95698 310874 95934
rect 310294 95614 310874 95698
rect 310294 95378 310466 95614
rect 310702 95378 310874 95614
rect 310294 59934 310874 95378
rect 310294 59698 310466 59934
rect 310702 59698 310874 59934
rect 310294 59614 310874 59698
rect 310294 59378 310466 59614
rect 310702 59378 310874 59614
rect 310294 23934 310874 59378
rect 310294 23698 310466 23934
rect 310702 23698 310874 23934
rect 310294 23614 310874 23698
rect 310294 23378 310466 23614
rect 310702 23378 310874 23614
rect 310294 -3106 310874 23378
rect 310294 -3342 310466 -3106
rect 310702 -3342 310874 -3106
rect 310294 -3426 310874 -3342
rect 310294 -3662 310466 -3426
rect 310702 -3662 310874 -3426
rect 310294 -3674 310874 -3662
rect 313774 675414 314354 708882
rect 313774 675178 313946 675414
rect 314182 675178 314354 675414
rect 313774 675094 314354 675178
rect 313774 674858 313946 675094
rect 314182 674858 314354 675094
rect 313774 639414 314354 674858
rect 313774 639178 313946 639414
rect 314182 639178 314354 639414
rect 313774 639094 314354 639178
rect 313774 638858 313946 639094
rect 314182 638858 314354 639094
rect 313774 603414 314354 638858
rect 313774 603178 313946 603414
rect 314182 603178 314354 603414
rect 313774 603094 314354 603178
rect 313774 602858 313946 603094
rect 314182 602858 314354 603094
rect 313774 567414 314354 602858
rect 313774 567178 313946 567414
rect 314182 567178 314354 567414
rect 313774 567094 314354 567178
rect 313774 566858 313946 567094
rect 314182 566858 314354 567094
rect 313774 531414 314354 566858
rect 313774 531178 313946 531414
rect 314182 531178 314354 531414
rect 313774 531094 314354 531178
rect 313774 530858 313946 531094
rect 314182 530858 314354 531094
rect 313774 495414 314354 530858
rect 313774 495178 313946 495414
rect 314182 495178 314354 495414
rect 313774 495094 314354 495178
rect 313774 494858 313946 495094
rect 314182 494858 314354 495094
rect 313774 459414 314354 494858
rect 313774 459178 313946 459414
rect 314182 459178 314354 459414
rect 313774 459094 314354 459178
rect 313774 458858 313946 459094
rect 314182 458858 314354 459094
rect 313774 423414 314354 458858
rect 313774 423178 313946 423414
rect 314182 423178 314354 423414
rect 313774 423094 314354 423178
rect 313774 422858 313946 423094
rect 314182 422858 314354 423094
rect 313774 387414 314354 422858
rect 313774 387178 313946 387414
rect 314182 387178 314354 387414
rect 313774 387094 314354 387178
rect 313774 386858 313946 387094
rect 314182 386858 314354 387094
rect 313774 351414 314354 386858
rect 313774 351178 313946 351414
rect 314182 351178 314354 351414
rect 313774 351094 314354 351178
rect 313774 350858 313946 351094
rect 314182 350858 314354 351094
rect 313774 315414 314354 350858
rect 313774 315178 313946 315414
rect 314182 315178 314354 315414
rect 313774 315094 314354 315178
rect 313774 314858 313946 315094
rect 314182 314858 314354 315094
rect 313774 279414 314354 314858
rect 313774 279178 313946 279414
rect 314182 279178 314354 279414
rect 313774 279094 314354 279178
rect 313774 278858 313946 279094
rect 314182 278858 314354 279094
rect 313774 243414 314354 278858
rect 313774 243178 313946 243414
rect 314182 243178 314354 243414
rect 313774 243094 314354 243178
rect 313774 242858 313946 243094
rect 314182 242858 314354 243094
rect 313774 207414 314354 242858
rect 313774 207178 313946 207414
rect 314182 207178 314354 207414
rect 313774 207094 314354 207178
rect 313774 206858 313946 207094
rect 314182 206858 314354 207094
rect 313774 171414 314354 206858
rect 313774 171178 313946 171414
rect 314182 171178 314354 171414
rect 313774 171094 314354 171178
rect 313774 170858 313946 171094
rect 314182 170858 314354 171094
rect 313774 135414 314354 170858
rect 313774 135178 313946 135414
rect 314182 135178 314354 135414
rect 313774 135094 314354 135178
rect 313774 134858 313946 135094
rect 314182 134858 314354 135094
rect 313774 99414 314354 134858
rect 313774 99178 313946 99414
rect 314182 99178 314354 99414
rect 313774 99094 314354 99178
rect 313774 98858 313946 99094
rect 314182 98858 314354 99094
rect 313774 63414 314354 98858
rect 313774 63178 313946 63414
rect 314182 63178 314354 63414
rect 313774 63094 314354 63178
rect 313774 62858 313946 63094
rect 314182 62858 314354 63094
rect 313774 27414 314354 62858
rect 313774 27178 313946 27414
rect 314182 27178 314354 27414
rect 313774 27094 314354 27178
rect 313774 26858 313946 27094
rect 314182 26858 314354 27094
rect 313774 -4946 314354 26858
rect 313774 -5182 313946 -4946
rect 314182 -5182 314354 -4946
rect 313774 -5266 314354 -5182
rect 313774 -5502 313946 -5266
rect 314182 -5502 314354 -5266
rect 313774 -5514 314354 -5502
rect 317254 678894 317834 710722
rect 335254 710358 335834 711290
rect 335254 710122 335426 710358
rect 335662 710122 335834 710358
rect 335254 710038 335834 710122
rect 335254 709802 335426 710038
rect 335662 709802 335834 710038
rect 331774 708518 332354 709450
rect 331774 708282 331946 708518
rect 332182 708282 332354 708518
rect 331774 708198 332354 708282
rect 331774 707962 331946 708198
rect 332182 707962 332354 708198
rect 328294 706678 328874 707610
rect 328294 706442 328466 706678
rect 328702 706442 328874 706678
rect 328294 706358 328874 706442
rect 328294 706122 328466 706358
rect 328702 706122 328874 706358
rect 317254 678658 317426 678894
rect 317662 678658 317834 678894
rect 317254 678574 317834 678658
rect 317254 678338 317426 678574
rect 317662 678338 317834 678574
rect 317254 642894 317834 678338
rect 317254 642658 317426 642894
rect 317662 642658 317834 642894
rect 317254 642574 317834 642658
rect 317254 642338 317426 642574
rect 317662 642338 317834 642574
rect 317254 606894 317834 642338
rect 317254 606658 317426 606894
rect 317662 606658 317834 606894
rect 317254 606574 317834 606658
rect 317254 606338 317426 606574
rect 317662 606338 317834 606574
rect 317254 570894 317834 606338
rect 317254 570658 317426 570894
rect 317662 570658 317834 570894
rect 317254 570574 317834 570658
rect 317254 570338 317426 570574
rect 317662 570338 317834 570574
rect 317254 534894 317834 570338
rect 317254 534658 317426 534894
rect 317662 534658 317834 534894
rect 317254 534574 317834 534658
rect 317254 534338 317426 534574
rect 317662 534338 317834 534574
rect 317254 498894 317834 534338
rect 317254 498658 317426 498894
rect 317662 498658 317834 498894
rect 317254 498574 317834 498658
rect 317254 498338 317426 498574
rect 317662 498338 317834 498574
rect 317254 462894 317834 498338
rect 317254 462658 317426 462894
rect 317662 462658 317834 462894
rect 317254 462574 317834 462658
rect 317254 462338 317426 462574
rect 317662 462338 317834 462574
rect 317254 426894 317834 462338
rect 317254 426658 317426 426894
rect 317662 426658 317834 426894
rect 317254 426574 317834 426658
rect 317254 426338 317426 426574
rect 317662 426338 317834 426574
rect 317254 390894 317834 426338
rect 317254 390658 317426 390894
rect 317662 390658 317834 390894
rect 317254 390574 317834 390658
rect 317254 390338 317426 390574
rect 317662 390338 317834 390574
rect 317254 354894 317834 390338
rect 317254 354658 317426 354894
rect 317662 354658 317834 354894
rect 317254 354574 317834 354658
rect 317254 354338 317426 354574
rect 317662 354338 317834 354574
rect 317254 318894 317834 354338
rect 317254 318658 317426 318894
rect 317662 318658 317834 318894
rect 317254 318574 317834 318658
rect 317254 318338 317426 318574
rect 317662 318338 317834 318574
rect 317254 282894 317834 318338
rect 317254 282658 317426 282894
rect 317662 282658 317834 282894
rect 317254 282574 317834 282658
rect 317254 282338 317426 282574
rect 317662 282338 317834 282574
rect 317254 246894 317834 282338
rect 317254 246658 317426 246894
rect 317662 246658 317834 246894
rect 317254 246574 317834 246658
rect 317254 246338 317426 246574
rect 317662 246338 317834 246574
rect 317254 210894 317834 246338
rect 317254 210658 317426 210894
rect 317662 210658 317834 210894
rect 317254 210574 317834 210658
rect 317254 210338 317426 210574
rect 317662 210338 317834 210574
rect 317254 174894 317834 210338
rect 317254 174658 317426 174894
rect 317662 174658 317834 174894
rect 317254 174574 317834 174658
rect 317254 174338 317426 174574
rect 317662 174338 317834 174574
rect 317254 138894 317834 174338
rect 317254 138658 317426 138894
rect 317662 138658 317834 138894
rect 317254 138574 317834 138658
rect 317254 138338 317426 138574
rect 317662 138338 317834 138574
rect 317254 102894 317834 138338
rect 317254 102658 317426 102894
rect 317662 102658 317834 102894
rect 317254 102574 317834 102658
rect 317254 102338 317426 102574
rect 317662 102338 317834 102574
rect 317254 66894 317834 102338
rect 317254 66658 317426 66894
rect 317662 66658 317834 66894
rect 317254 66574 317834 66658
rect 317254 66338 317426 66574
rect 317662 66338 317834 66574
rect 317254 30894 317834 66338
rect 317254 30658 317426 30894
rect 317662 30658 317834 30894
rect 317254 30574 317834 30658
rect 317254 30338 317426 30574
rect 317662 30338 317834 30574
rect 299254 -6102 299426 -5866
rect 299662 -6102 299834 -5866
rect 299254 -6186 299834 -6102
rect 299254 -6422 299426 -6186
rect 299662 -6422 299834 -6186
rect 299254 -7354 299834 -6422
rect 317254 -6786 317834 30338
rect 324814 704838 325394 705770
rect 324814 704602 324986 704838
rect 325222 704602 325394 704838
rect 324814 704518 325394 704602
rect 324814 704282 324986 704518
rect 325222 704282 325394 704518
rect 324814 686454 325394 704282
rect 324814 686218 324986 686454
rect 325222 686218 325394 686454
rect 324814 686134 325394 686218
rect 324814 685898 324986 686134
rect 325222 685898 325394 686134
rect 324814 650454 325394 685898
rect 324814 650218 324986 650454
rect 325222 650218 325394 650454
rect 324814 650134 325394 650218
rect 324814 649898 324986 650134
rect 325222 649898 325394 650134
rect 324814 614454 325394 649898
rect 324814 614218 324986 614454
rect 325222 614218 325394 614454
rect 324814 614134 325394 614218
rect 324814 613898 324986 614134
rect 325222 613898 325394 614134
rect 324814 578454 325394 613898
rect 324814 578218 324986 578454
rect 325222 578218 325394 578454
rect 324814 578134 325394 578218
rect 324814 577898 324986 578134
rect 325222 577898 325394 578134
rect 324814 542454 325394 577898
rect 324814 542218 324986 542454
rect 325222 542218 325394 542454
rect 324814 542134 325394 542218
rect 324814 541898 324986 542134
rect 325222 541898 325394 542134
rect 324814 506454 325394 541898
rect 324814 506218 324986 506454
rect 325222 506218 325394 506454
rect 324814 506134 325394 506218
rect 324814 505898 324986 506134
rect 325222 505898 325394 506134
rect 324814 470454 325394 505898
rect 324814 470218 324986 470454
rect 325222 470218 325394 470454
rect 324814 470134 325394 470218
rect 324814 469898 324986 470134
rect 325222 469898 325394 470134
rect 324814 434454 325394 469898
rect 324814 434218 324986 434454
rect 325222 434218 325394 434454
rect 324814 434134 325394 434218
rect 324814 433898 324986 434134
rect 325222 433898 325394 434134
rect 324814 398454 325394 433898
rect 324814 398218 324986 398454
rect 325222 398218 325394 398454
rect 324814 398134 325394 398218
rect 324814 397898 324986 398134
rect 325222 397898 325394 398134
rect 324814 362454 325394 397898
rect 324814 362218 324986 362454
rect 325222 362218 325394 362454
rect 324814 362134 325394 362218
rect 324814 361898 324986 362134
rect 325222 361898 325394 362134
rect 324814 326454 325394 361898
rect 324814 326218 324986 326454
rect 325222 326218 325394 326454
rect 324814 326134 325394 326218
rect 324814 325898 324986 326134
rect 325222 325898 325394 326134
rect 324814 290454 325394 325898
rect 324814 290218 324986 290454
rect 325222 290218 325394 290454
rect 324814 290134 325394 290218
rect 324814 289898 324986 290134
rect 325222 289898 325394 290134
rect 324814 254454 325394 289898
rect 324814 254218 324986 254454
rect 325222 254218 325394 254454
rect 324814 254134 325394 254218
rect 324814 253898 324986 254134
rect 325222 253898 325394 254134
rect 324814 218454 325394 253898
rect 324814 218218 324986 218454
rect 325222 218218 325394 218454
rect 324814 218134 325394 218218
rect 324814 217898 324986 218134
rect 325222 217898 325394 218134
rect 324814 182454 325394 217898
rect 324814 182218 324986 182454
rect 325222 182218 325394 182454
rect 324814 182134 325394 182218
rect 324814 181898 324986 182134
rect 325222 181898 325394 182134
rect 324814 146454 325394 181898
rect 324814 146218 324986 146454
rect 325222 146218 325394 146454
rect 324814 146134 325394 146218
rect 324814 145898 324986 146134
rect 325222 145898 325394 146134
rect 324814 110454 325394 145898
rect 324814 110218 324986 110454
rect 325222 110218 325394 110454
rect 324814 110134 325394 110218
rect 324814 109898 324986 110134
rect 325222 109898 325394 110134
rect 324814 74454 325394 109898
rect 324814 74218 324986 74454
rect 325222 74218 325394 74454
rect 324814 74134 325394 74218
rect 324814 73898 324986 74134
rect 325222 73898 325394 74134
rect 324814 38454 325394 73898
rect 324814 38218 324986 38454
rect 325222 38218 325394 38454
rect 324814 38134 325394 38218
rect 324814 37898 324986 38134
rect 325222 37898 325394 38134
rect 324814 2454 325394 37898
rect 324814 2218 324986 2454
rect 325222 2218 325394 2454
rect 324814 2134 325394 2218
rect 324814 1898 324986 2134
rect 325222 1898 325394 2134
rect 324814 -346 325394 1898
rect 324814 -582 324986 -346
rect 325222 -582 325394 -346
rect 324814 -666 325394 -582
rect 324814 -902 324986 -666
rect 325222 -902 325394 -666
rect 324814 -1834 325394 -902
rect 328294 689934 328874 706122
rect 328294 689698 328466 689934
rect 328702 689698 328874 689934
rect 328294 689614 328874 689698
rect 328294 689378 328466 689614
rect 328702 689378 328874 689614
rect 328294 653934 328874 689378
rect 328294 653698 328466 653934
rect 328702 653698 328874 653934
rect 328294 653614 328874 653698
rect 328294 653378 328466 653614
rect 328702 653378 328874 653614
rect 328294 617934 328874 653378
rect 328294 617698 328466 617934
rect 328702 617698 328874 617934
rect 328294 617614 328874 617698
rect 328294 617378 328466 617614
rect 328702 617378 328874 617614
rect 328294 581934 328874 617378
rect 328294 581698 328466 581934
rect 328702 581698 328874 581934
rect 328294 581614 328874 581698
rect 328294 581378 328466 581614
rect 328702 581378 328874 581614
rect 328294 545934 328874 581378
rect 328294 545698 328466 545934
rect 328702 545698 328874 545934
rect 328294 545614 328874 545698
rect 328294 545378 328466 545614
rect 328702 545378 328874 545614
rect 328294 509934 328874 545378
rect 328294 509698 328466 509934
rect 328702 509698 328874 509934
rect 328294 509614 328874 509698
rect 328294 509378 328466 509614
rect 328702 509378 328874 509614
rect 328294 473934 328874 509378
rect 328294 473698 328466 473934
rect 328702 473698 328874 473934
rect 328294 473614 328874 473698
rect 328294 473378 328466 473614
rect 328702 473378 328874 473614
rect 328294 437934 328874 473378
rect 328294 437698 328466 437934
rect 328702 437698 328874 437934
rect 328294 437614 328874 437698
rect 328294 437378 328466 437614
rect 328702 437378 328874 437614
rect 328294 401934 328874 437378
rect 328294 401698 328466 401934
rect 328702 401698 328874 401934
rect 328294 401614 328874 401698
rect 328294 401378 328466 401614
rect 328702 401378 328874 401614
rect 328294 365934 328874 401378
rect 328294 365698 328466 365934
rect 328702 365698 328874 365934
rect 328294 365614 328874 365698
rect 328294 365378 328466 365614
rect 328702 365378 328874 365614
rect 328294 329934 328874 365378
rect 328294 329698 328466 329934
rect 328702 329698 328874 329934
rect 328294 329614 328874 329698
rect 328294 329378 328466 329614
rect 328702 329378 328874 329614
rect 328294 293934 328874 329378
rect 328294 293698 328466 293934
rect 328702 293698 328874 293934
rect 328294 293614 328874 293698
rect 328294 293378 328466 293614
rect 328702 293378 328874 293614
rect 328294 257934 328874 293378
rect 328294 257698 328466 257934
rect 328702 257698 328874 257934
rect 328294 257614 328874 257698
rect 328294 257378 328466 257614
rect 328702 257378 328874 257614
rect 328294 221934 328874 257378
rect 328294 221698 328466 221934
rect 328702 221698 328874 221934
rect 328294 221614 328874 221698
rect 328294 221378 328466 221614
rect 328702 221378 328874 221614
rect 328294 185934 328874 221378
rect 328294 185698 328466 185934
rect 328702 185698 328874 185934
rect 328294 185614 328874 185698
rect 328294 185378 328466 185614
rect 328702 185378 328874 185614
rect 328294 149934 328874 185378
rect 328294 149698 328466 149934
rect 328702 149698 328874 149934
rect 328294 149614 328874 149698
rect 328294 149378 328466 149614
rect 328702 149378 328874 149614
rect 328294 113934 328874 149378
rect 328294 113698 328466 113934
rect 328702 113698 328874 113934
rect 328294 113614 328874 113698
rect 328294 113378 328466 113614
rect 328702 113378 328874 113614
rect 328294 77934 328874 113378
rect 328294 77698 328466 77934
rect 328702 77698 328874 77934
rect 328294 77614 328874 77698
rect 328294 77378 328466 77614
rect 328702 77378 328874 77614
rect 328294 41934 328874 77378
rect 328294 41698 328466 41934
rect 328702 41698 328874 41934
rect 328294 41614 328874 41698
rect 328294 41378 328466 41614
rect 328702 41378 328874 41614
rect 328294 5934 328874 41378
rect 328294 5698 328466 5934
rect 328702 5698 328874 5934
rect 328294 5614 328874 5698
rect 328294 5378 328466 5614
rect 328702 5378 328874 5614
rect 328294 -2186 328874 5378
rect 328294 -2422 328466 -2186
rect 328702 -2422 328874 -2186
rect 328294 -2506 328874 -2422
rect 328294 -2742 328466 -2506
rect 328702 -2742 328874 -2506
rect 328294 -3674 328874 -2742
rect 331774 693414 332354 707962
rect 331774 693178 331946 693414
rect 332182 693178 332354 693414
rect 331774 693094 332354 693178
rect 331774 692858 331946 693094
rect 332182 692858 332354 693094
rect 331774 657414 332354 692858
rect 331774 657178 331946 657414
rect 332182 657178 332354 657414
rect 331774 657094 332354 657178
rect 331774 656858 331946 657094
rect 332182 656858 332354 657094
rect 331774 621414 332354 656858
rect 331774 621178 331946 621414
rect 332182 621178 332354 621414
rect 331774 621094 332354 621178
rect 331774 620858 331946 621094
rect 332182 620858 332354 621094
rect 331774 585414 332354 620858
rect 331774 585178 331946 585414
rect 332182 585178 332354 585414
rect 331774 585094 332354 585178
rect 331774 584858 331946 585094
rect 332182 584858 332354 585094
rect 331774 549414 332354 584858
rect 331774 549178 331946 549414
rect 332182 549178 332354 549414
rect 331774 549094 332354 549178
rect 331774 548858 331946 549094
rect 332182 548858 332354 549094
rect 331774 513414 332354 548858
rect 331774 513178 331946 513414
rect 332182 513178 332354 513414
rect 331774 513094 332354 513178
rect 331774 512858 331946 513094
rect 332182 512858 332354 513094
rect 331774 477414 332354 512858
rect 331774 477178 331946 477414
rect 332182 477178 332354 477414
rect 331774 477094 332354 477178
rect 331774 476858 331946 477094
rect 332182 476858 332354 477094
rect 331774 441414 332354 476858
rect 331774 441178 331946 441414
rect 332182 441178 332354 441414
rect 331774 441094 332354 441178
rect 331774 440858 331946 441094
rect 332182 440858 332354 441094
rect 331774 405414 332354 440858
rect 331774 405178 331946 405414
rect 332182 405178 332354 405414
rect 331774 405094 332354 405178
rect 331774 404858 331946 405094
rect 332182 404858 332354 405094
rect 331774 369414 332354 404858
rect 331774 369178 331946 369414
rect 332182 369178 332354 369414
rect 331774 369094 332354 369178
rect 331774 368858 331946 369094
rect 332182 368858 332354 369094
rect 331774 333414 332354 368858
rect 331774 333178 331946 333414
rect 332182 333178 332354 333414
rect 331774 333094 332354 333178
rect 331774 332858 331946 333094
rect 332182 332858 332354 333094
rect 331774 297414 332354 332858
rect 331774 297178 331946 297414
rect 332182 297178 332354 297414
rect 331774 297094 332354 297178
rect 331774 296858 331946 297094
rect 332182 296858 332354 297094
rect 331774 261414 332354 296858
rect 331774 261178 331946 261414
rect 332182 261178 332354 261414
rect 331774 261094 332354 261178
rect 331774 260858 331946 261094
rect 332182 260858 332354 261094
rect 331774 225414 332354 260858
rect 331774 225178 331946 225414
rect 332182 225178 332354 225414
rect 331774 225094 332354 225178
rect 331774 224858 331946 225094
rect 332182 224858 332354 225094
rect 331774 189414 332354 224858
rect 331774 189178 331946 189414
rect 332182 189178 332354 189414
rect 331774 189094 332354 189178
rect 331774 188858 331946 189094
rect 332182 188858 332354 189094
rect 331774 153414 332354 188858
rect 331774 153178 331946 153414
rect 332182 153178 332354 153414
rect 331774 153094 332354 153178
rect 331774 152858 331946 153094
rect 332182 152858 332354 153094
rect 331774 117414 332354 152858
rect 331774 117178 331946 117414
rect 332182 117178 332354 117414
rect 331774 117094 332354 117178
rect 331774 116858 331946 117094
rect 332182 116858 332354 117094
rect 331774 81414 332354 116858
rect 331774 81178 331946 81414
rect 332182 81178 332354 81414
rect 331774 81094 332354 81178
rect 331774 80858 331946 81094
rect 332182 80858 332354 81094
rect 331774 45414 332354 80858
rect 331774 45178 331946 45414
rect 332182 45178 332354 45414
rect 331774 45094 332354 45178
rect 331774 44858 331946 45094
rect 332182 44858 332354 45094
rect 331774 9414 332354 44858
rect 331774 9178 331946 9414
rect 332182 9178 332354 9414
rect 331774 9094 332354 9178
rect 331774 8858 331946 9094
rect 332182 8858 332354 9094
rect 331774 -4026 332354 8858
rect 331774 -4262 331946 -4026
rect 332182 -4262 332354 -4026
rect 331774 -4346 332354 -4262
rect 331774 -4582 331946 -4346
rect 332182 -4582 332354 -4346
rect 331774 -5514 332354 -4582
rect 335254 696894 335834 709802
rect 353254 711278 353834 711290
rect 353254 711042 353426 711278
rect 353662 711042 353834 711278
rect 353254 710958 353834 711042
rect 353254 710722 353426 710958
rect 353662 710722 353834 710958
rect 349774 709438 350354 709450
rect 349774 709202 349946 709438
rect 350182 709202 350354 709438
rect 349774 709118 350354 709202
rect 349774 708882 349946 709118
rect 350182 708882 350354 709118
rect 346294 707598 346874 707610
rect 346294 707362 346466 707598
rect 346702 707362 346874 707598
rect 346294 707278 346874 707362
rect 346294 707042 346466 707278
rect 346702 707042 346874 707278
rect 335254 696658 335426 696894
rect 335662 696658 335834 696894
rect 335254 696574 335834 696658
rect 335254 696338 335426 696574
rect 335662 696338 335834 696574
rect 335254 660894 335834 696338
rect 335254 660658 335426 660894
rect 335662 660658 335834 660894
rect 335254 660574 335834 660658
rect 335254 660338 335426 660574
rect 335662 660338 335834 660574
rect 335254 624894 335834 660338
rect 335254 624658 335426 624894
rect 335662 624658 335834 624894
rect 335254 624574 335834 624658
rect 335254 624338 335426 624574
rect 335662 624338 335834 624574
rect 335254 588894 335834 624338
rect 335254 588658 335426 588894
rect 335662 588658 335834 588894
rect 335254 588574 335834 588658
rect 335254 588338 335426 588574
rect 335662 588338 335834 588574
rect 335254 552894 335834 588338
rect 335254 552658 335426 552894
rect 335662 552658 335834 552894
rect 335254 552574 335834 552658
rect 335254 552338 335426 552574
rect 335662 552338 335834 552574
rect 335254 516894 335834 552338
rect 335254 516658 335426 516894
rect 335662 516658 335834 516894
rect 335254 516574 335834 516658
rect 335254 516338 335426 516574
rect 335662 516338 335834 516574
rect 335254 480894 335834 516338
rect 335254 480658 335426 480894
rect 335662 480658 335834 480894
rect 335254 480574 335834 480658
rect 335254 480338 335426 480574
rect 335662 480338 335834 480574
rect 335254 444894 335834 480338
rect 335254 444658 335426 444894
rect 335662 444658 335834 444894
rect 335254 444574 335834 444658
rect 335254 444338 335426 444574
rect 335662 444338 335834 444574
rect 335254 408894 335834 444338
rect 335254 408658 335426 408894
rect 335662 408658 335834 408894
rect 335254 408574 335834 408658
rect 335254 408338 335426 408574
rect 335662 408338 335834 408574
rect 335254 372894 335834 408338
rect 335254 372658 335426 372894
rect 335662 372658 335834 372894
rect 335254 372574 335834 372658
rect 335254 372338 335426 372574
rect 335662 372338 335834 372574
rect 335254 336894 335834 372338
rect 335254 336658 335426 336894
rect 335662 336658 335834 336894
rect 335254 336574 335834 336658
rect 335254 336338 335426 336574
rect 335662 336338 335834 336574
rect 335254 300894 335834 336338
rect 335254 300658 335426 300894
rect 335662 300658 335834 300894
rect 335254 300574 335834 300658
rect 335254 300338 335426 300574
rect 335662 300338 335834 300574
rect 335254 264894 335834 300338
rect 335254 264658 335426 264894
rect 335662 264658 335834 264894
rect 335254 264574 335834 264658
rect 335254 264338 335426 264574
rect 335662 264338 335834 264574
rect 335254 228894 335834 264338
rect 335254 228658 335426 228894
rect 335662 228658 335834 228894
rect 335254 228574 335834 228658
rect 335254 228338 335426 228574
rect 335662 228338 335834 228574
rect 335254 192894 335834 228338
rect 335254 192658 335426 192894
rect 335662 192658 335834 192894
rect 335254 192574 335834 192658
rect 335254 192338 335426 192574
rect 335662 192338 335834 192574
rect 335254 156894 335834 192338
rect 335254 156658 335426 156894
rect 335662 156658 335834 156894
rect 335254 156574 335834 156658
rect 335254 156338 335426 156574
rect 335662 156338 335834 156574
rect 335254 120894 335834 156338
rect 335254 120658 335426 120894
rect 335662 120658 335834 120894
rect 335254 120574 335834 120658
rect 335254 120338 335426 120574
rect 335662 120338 335834 120574
rect 335254 84894 335834 120338
rect 335254 84658 335426 84894
rect 335662 84658 335834 84894
rect 335254 84574 335834 84658
rect 335254 84338 335426 84574
rect 335662 84338 335834 84574
rect 335254 48894 335834 84338
rect 335254 48658 335426 48894
rect 335662 48658 335834 48894
rect 335254 48574 335834 48658
rect 335254 48338 335426 48574
rect 335662 48338 335834 48574
rect 335254 12894 335834 48338
rect 335254 12658 335426 12894
rect 335662 12658 335834 12894
rect 335254 12574 335834 12658
rect 335254 12338 335426 12574
rect 335662 12338 335834 12574
rect 317254 -7022 317426 -6786
rect 317662 -7022 317834 -6786
rect 317254 -7106 317834 -7022
rect 317254 -7342 317426 -7106
rect 317662 -7342 317834 -7106
rect 317254 -7354 317834 -7342
rect 335254 -5866 335834 12338
rect 342814 705758 343394 705770
rect 342814 705522 342986 705758
rect 343222 705522 343394 705758
rect 342814 705438 343394 705522
rect 342814 705202 342986 705438
rect 343222 705202 343394 705438
rect 342814 668454 343394 705202
rect 342814 668218 342986 668454
rect 343222 668218 343394 668454
rect 342814 668134 343394 668218
rect 342814 667898 342986 668134
rect 343222 667898 343394 668134
rect 342814 632454 343394 667898
rect 342814 632218 342986 632454
rect 343222 632218 343394 632454
rect 342814 632134 343394 632218
rect 342814 631898 342986 632134
rect 343222 631898 343394 632134
rect 342814 596454 343394 631898
rect 342814 596218 342986 596454
rect 343222 596218 343394 596454
rect 342814 596134 343394 596218
rect 342814 595898 342986 596134
rect 343222 595898 343394 596134
rect 342814 560454 343394 595898
rect 342814 560218 342986 560454
rect 343222 560218 343394 560454
rect 342814 560134 343394 560218
rect 342814 559898 342986 560134
rect 343222 559898 343394 560134
rect 342814 524454 343394 559898
rect 342814 524218 342986 524454
rect 343222 524218 343394 524454
rect 342814 524134 343394 524218
rect 342814 523898 342986 524134
rect 343222 523898 343394 524134
rect 342814 488454 343394 523898
rect 342814 488218 342986 488454
rect 343222 488218 343394 488454
rect 342814 488134 343394 488218
rect 342814 487898 342986 488134
rect 343222 487898 343394 488134
rect 342814 452454 343394 487898
rect 342814 452218 342986 452454
rect 343222 452218 343394 452454
rect 342814 452134 343394 452218
rect 342814 451898 342986 452134
rect 343222 451898 343394 452134
rect 342814 416454 343394 451898
rect 342814 416218 342986 416454
rect 343222 416218 343394 416454
rect 342814 416134 343394 416218
rect 342814 415898 342986 416134
rect 343222 415898 343394 416134
rect 342814 380454 343394 415898
rect 342814 380218 342986 380454
rect 343222 380218 343394 380454
rect 342814 380134 343394 380218
rect 342814 379898 342986 380134
rect 343222 379898 343394 380134
rect 342814 344454 343394 379898
rect 346294 671934 346874 707042
rect 346294 671698 346466 671934
rect 346702 671698 346874 671934
rect 346294 671614 346874 671698
rect 346294 671378 346466 671614
rect 346702 671378 346874 671614
rect 346294 635934 346874 671378
rect 346294 635698 346466 635934
rect 346702 635698 346874 635934
rect 346294 635614 346874 635698
rect 346294 635378 346466 635614
rect 346702 635378 346874 635614
rect 346294 599934 346874 635378
rect 346294 599698 346466 599934
rect 346702 599698 346874 599934
rect 346294 599614 346874 599698
rect 346294 599378 346466 599614
rect 346702 599378 346874 599614
rect 346294 563934 346874 599378
rect 346294 563698 346466 563934
rect 346702 563698 346874 563934
rect 346294 563614 346874 563698
rect 346294 563378 346466 563614
rect 346702 563378 346874 563614
rect 346294 527934 346874 563378
rect 346294 527698 346466 527934
rect 346702 527698 346874 527934
rect 346294 527614 346874 527698
rect 346294 527378 346466 527614
rect 346702 527378 346874 527614
rect 346294 491934 346874 527378
rect 346294 491698 346466 491934
rect 346702 491698 346874 491934
rect 346294 491614 346874 491698
rect 346294 491378 346466 491614
rect 346702 491378 346874 491614
rect 346294 455934 346874 491378
rect 346294 455698 346466 455934
rect 346702 455698 346874 455934
rect 346294 455614 346874 455698
rect 346294 455378 346466 455614
rect 346702 455378 346874 455614
rect 346294 419934 346874 455378
rect 346294 419698 346466 419934
rect 346702 419698 346874 419934
rect 346294 419614 346874 419698
rect 346294 419378 346466 419614
rect 346702 419378 346874 419614
rect 346294 383934 346874 419378
rect 346294 383698 346466 383934
rect 346702 383698 346874 383934
rect 346294 383614 346874 383698
rect 346294 383378 346466 383614
rect 346702 383378 346874 383614
rect 344878 360858 344938 363342
rect 342814 344218 342986 344454
rect 343222 344218 343394 344454
rect 342814 344134 343394 344218
rect 342814 343898 342986 344134
rect 343222 343898 343394 344134
rect 342814 308454 343394 343898
rect 342814 308218 342986 308454
rect 343222 308218 343394 308454
rect 342814 308134 343394 308218
rect 342814 307898 342986 308134
rect 343222 307898 343394 308134
rect 342814 272454 343394 307898
rect 342814 272218 342986 272454
rect 343222 272218 343394 272454
rect 342814 272134 343394 272218
rect 342814 271898 342986 272134
rect 343222 271898 343394 272134
rect 342814 236454 343394 271898
rect 342814 236218 342986 236454
rect 343222 236218 343394 236454
rect 342814 236134 343394 236218
rect 342814 235898 342986 236134
rect 343222 235898 343394 236134
rect 342814 200454 343394 235898
rect 342814 200218 342986 200454
rect 343222 200218 343394 200454
rect 342814 200134 343394 200218
rect 342814 199898 342986 200134
rect 343222 199898 343394 200134
rect 342814 164454 343394 199898
rect 342814 164218 342986 164454
rect 343222 164218 343394 164454
rect 342814 164134 343394 164218
rect 342814 163898 342986 164134
rect 343222 163898 343394 164134
rect 342814 128454 343394 163898
rect 342814 128218 342986 128454
rect 343222 128218 343394 128454
rect 342814 128134 343394 128218
rect 342814 127898 342986 128134
rect 343222 127898 343394 128134
rect 342814 92454 343394 127898
rect 342814 92218 342986 92454
rect 343222 92218 343394 92454
rect 342814 92134 343394 92218
rect 342814 91898 342986 92134
rect 343222 91898 343394 92134
rect 342814 56454 343394 91898
rect 342814 56218 342986 56454
rect 343222 56218 343394 56454
rect 342814 56134 343394 56218
rect 342814 55898 342986 56134
rect 343222 55898 343394 56134
rect 342814 20454 343394 55898
rect 342814 20218 342986 20454
rect 343222 20218 343394 20454
rect 342814 20134 343394 20218
rect 342814 19898 342986 20134
rect 343222 19898 343394 20134
rect 342814 -1266 343394 19898
rect 342814 -1502 342986 -1266
rect 343222 -1502 343394 -1266
rect 342814 -1586 343394 -1502
rect 342814 -1822 342986 -1586
rect 343222 -1822 343394 -1586
rect 342814 -1834 343394 -1822
rect 346294 347934 346874 383378
rect 346294 347698 346466 347934
rect 346702 347698 346874 347934
rect 346294 347614 346874 347698
rect 346294 347378 346466 347614
rect 346702 347378 346874 347614
rect 346294 311934 346874 347378
rect 346294 311698 346466 311934
rect 346702 311698 346874 311934
rect 346294 311614 346874 311698
rect 346294 311378 346466 311614
rect 346702 311378 346874 311614
rect 346294 275934 346874 311378
rect 346294 275698 346466 275934
rect 346702 275698 346874 275934
rect 346294 275614 346874 275698
rect 346294 275378 346466 275614
rect 346702 275378 346874 275614
rect 346294 239934 346874 275378
rect 346294 239698 346466 239934
rect 346702 239698 346874 239934
rect 346294 239614 346874 239698
rect 346294 239378 346466 239614
rect 346702 239378 346874 239614
rect 346294 203934 346874 239378
rect 346294 203698 346466 203934
rect 346702 203698 346874 203934
rect 346294 203614 346874 203698
rect 346294 203378 346466 203614
rect 346702 203378 346874 203614
rect 346294 167934 346874 203378
rect 346294 167698 346466 167934
rect 346702 167698 346874 167934
rect 346294 167614 346874 167698
rect 346294 167378 346466 167614
rect 346702 167378 346874 167614
rect 346294 131934 346874 167378
rect 346294 131698 346466 131934
rect 346702 131698 346874 131934
rect 346294 131614 346874 131698
rect 346294 131378 346466 131614
rect 346702 131378 346874 131614
rect 346294 95934 346874 131378
rect 346294 95698 346466 95934
rect 346702 95698 346874 95934
rect 346294 95614 346874 95698
rect 346294 95378 346466 95614
rect 346702 95378 346874 95614
rect 346294 59934 346874 95378
rect 346294 59698 346466 59934
rect 346702 59698 346874 59934
rect 346294 59614 346874 59698
rect 346294 59378 346466 59614
rect 346702 59378 346874 59614
rect 346294 23934 346874 59378
rect 346294 23698 346466 23934
rect 346702 23698 346874 23934
rect 346294 23614 346874 23698
rect 346294 23378 346466 23614
rect 346702 23378 346874 23614
rect 346294 -3106 346874 23378
rect 346294 -3342 346466 -3106
rect 346702 -3342 346874 -3106
rect 346294 -3426 346874 -3342
rect 346294 -3662 346466 -3426
rect 346702 -3662 346874 -3426
rect 346294 -3674 346874 -3662
rect 349774 675414 350354 708882
rect 349774 675178 349946 675414
rect 350182 675178 350354 675414
rect 349774 675094 350354 675178
rect 349774 674858 349946 675094
rect 350182 674858 350354 675094
rect 349774 639414 350354 674858
rect 349774 639178 349946 639414
rect 350182 639178 350354 639414
rect 349774 639094 350354 639178
rect 349774 638858 349946 639094
rect 350182 638858 350354 639094
rect 349774 603414 350354 638858
rect 349774 603178 349946 603414
rect 350182 603178 350354 603414
rect 349774 603094 350354 603178
rect 349774 602858 349946 603094
rect 350182 602858 350354 603094
rect 349774 567414 350354 602858
rect 349774 567178 349946 567414
rect 350182 567178 350354 567414
rect 349774 567094 350354 567178
rect 349774 566858 349946 567094
rect 350182 566858 350354 567094
rect 349774 531414 350354 566858
rect 349774 531178 349946 531414
rect 350182 531178 350354 531414
rect 349774 531094 350354 531178
rect 349774 530858 349946 531094
rect 350182 530858 350354 531094
rect 349774 495414 350354 530858
rect 349774 495178 349946 495414
rect 350182 495178 350354 495414
rect 349774 495094 350354 495178
rect 349774 494858 349946 495094
rect 350182 494858 350354 495094
rect 349774 459414 350354 494858
rect 349774 459178 349946 459414
rect 350182 459178 350354 459414
rect 349774 459094 350354 459178
rect 349774 458858 349946 459094
rect 350182 458858 350354 459094
rect 349774 423414 350354 458858
rect 349774 423178 349946 423414
rect 350182 423178 350354 423414
rect 349774 423094 350354 423178
rect 349774 422858 349946 423094
rect 350182 422858 350354 423094
rect 349774 387414 350354 422858
rect 349774 387178 349946 387414
rect 350182 387178 350354 387414
rect 349774 387094 350354 387178
rect 349774 386858 349946 387094
rect 350182 386858 350354 387094
rect 349774 351414 350354 386858
rect 349774 351178 349946 351414
rect 350182 351178 350354 351414
rect 349774 351094 350354 351178
rect 349774 350858 349946 351094
rect 350182 350858 350354 351094
rect 349774 315414 350354 350858
rect 349774 315178 349946 315414
rect 350182 315178 350354 315414
rect 349774 315094 350354 315178
rect 349774 314858 349946 315094
rect 350182 314858 350354 315094
rect 349774 279414 350354 314858
rect 349774 279178 349946 279414
rect 350182 279178 350354 279414
rect 349774 279094 350354 279178
rect 349774 278858 349946 279094
rect 350182 278858 350354 279094
rect 349774 243414 350354 278858
rect 349774 243178 349946 243414
rect 350182 243178 350354 243414
rect 349774 243094 350354 243178
rect 349774 242858 349946 243094
rect 350182 242858 350354 243094
rect 349774 207414 350354 242858
rect 349774 207178 349946 207414
rect 350182 207178 350354 207414
rect 349774 207094 350354 207178
rect 349774 206858 349946 207094
rect 350182 206858 350354 207094
rect 349774 171414 350354 206858
rect 349774 171178 349946 171414
rect 350182 171178 350354 171414
rect 349774 171094 350354 171178
rect 349774 170858 349946 171094
rect 350182 170858 350354 171094
rect 349774 135414 350354 170858
rect 349774 135178 349946 135414
rect 350182 135178 350354 135414
rect 349774 135094 350354 135178
rect 349774 134858 349946 135094
rect 350182 134858 350354 135094
rect 349774 99414 350354 134858
rect 349774 99178 349946 99414
rect 350182 99178 350354 99414
rect 349774 99094 350354 99178
rect 349774 98858 349946 99094
rect 350182 98858 350354 99094
rect 349774 63414 350354 98858
rect 349774 63178 349946 63414
rect 350182 63178 350354 63414
rect 349774 63094 350354 63178
rect 349774 62858 349946 63094
rect 350182 62858 350354 63094
rect 349774 27414 350354 62858
rect 349774 27178 349946 27414
rect 350182 27178 350354 27414
rect 349774 27094 350354 27178
rect 349774 26858 349946 27094
rect 350182 26858 350354 27094
rect 349774 -4946 350354 26858
rect 349774 -5182 349946 -4946
rect 350182 -5182 350354 -4946
rect 349774 -5266 350354 -5182
rect 349774 -5502 349946 -5266
rect 350182 -5502 350354 -5266
rect 349774 -5514 350354 -5502
rect 353254 678894 353834 710722
rect 371254 710358 371834 711290
rect 371254 710122 371426 710358
rect 371662 710122 371834 710358
rect 371254 710038 371834 710122
rect 371254 709802 371426 710038
rect 371662 709802 371834 710038
rect 367774 708518 368354 709450
rect 367774 708282 367946 708518
rect 368182 708282 368354 708518
rect 367774 708198 368354 708282
rect 367774 707962 367946 708198
rect 368182 707962 368354 708198
rect 364294 706678 364874 707610
rect 364294 706442 364466 706678
rect 364702 706442 364874 706678
rect 364294 706358 364874 706442
rect 364294 706122 364466 706358
rect 364702 706122 364874 706358
rect 353254 678658 353426 678894
rect 353662 678658 353834 678894
rect 353254 678574 353834 678658
rect 353254 678338 353426 678574
rect 353662 678338 353834 678574
rect 353254 642894 353834 678338
rect 353254 642658 353426 642894
rect 353662 642658 353834 642894
rect 353254 642574 353834 642658
rect 353254 642338 353426 642574
rect 353662 642338 353834 642574
rect 353254 606894 353834 642338
rect 353254 606658 353426 606894
rect 353662 606658 353834 606894
rect 353254 606574 353834 606658
rect 353254 606338 353426 606574
rect 353662 606338 353834 606574
rect 353254 570894 353834 606338
rect 353254 570658 353426 570894
rect 353662 570658 353834 570894
rect 353254 570574 353834 570658
rect 353254 570338 353426 570574
rect 353662 570338 353834 570574
rect 353254 534894 353834 570338
rect 353254 534658 353426 534894
rect 353662 534658 353834 534894
rect 353254 534574 353834 534658
rect 353254 534338 353426 534574
rect 353662 534338 353834 534574
rect 353254 498894 353834 534338
rect 353254 498658 353426 498894
rect 353662 498658 353834 498894
rect 353254 498574 353834 498658
rect 353254 498338 353426 498574
rect 353662 498338 353834 498574
rect 353254 462894 353834 498338
rect 353254 462658 353426 462894
rect 353662 462658 353834 462894
rect 353254 462574 353834 462658
rect 353254 462338 353426 462574
rect 353662 462338 353834 462574
rect 353254 426894 353834 462338
rect 353254 426658 353426 426894
rect 353662 426658 353834 426894
rect 353254 426574 353834 426658
rect 353254 426338 353426 426574
rect 353662 426338 353834 426574
rect 353254 390894 353834 426338
rect 353254 390658 353426 390894
rect 353662 390658 353834 390894
rect 353254 390574 353834 390658
rect 353254 390338 353426 390574
rect 353662 390338 353834 390574
rect 353254 354894 353834 390338
rect 360814 704838 361394 705770
rect 360814 704602 360986 704838
rect 361222 704602 361394 704838
rect 360814 704518 361394 704602
rect 360814 704282 360986 704518
rect 361222 704282 361394 704518
rect 360814 686454 361394 704282
rect 360814 686218 360986 686454
rect 361222 686218 361394 686454
rect 360814 686134 361394 686218
rect 360814 685898 360986 686134
rect 361222 685898 361394 686134
rect 360814 650454 361394 685898
rect 360814 650218 360986 650454
rect 361222 650218 361394 650454
rect 360814 650134 361394 650218
rect 360814 649898 360986 650134
rect 361222 649898 361394 650134
rect 360814 614454 361394 649898
rect 360814 614218 360986 614454
rect 361222 614218 361394 614454
rect 360814 614134 361394 614218
rect 360814 613898 360986 614134
rect 361222 613898 361394 614134
rect 360814 578454 361394 613898
rect 360814 578218 360986 578454
rect 361222 578218 361394 578454
rect 360814 578134 361394 578218
rect 360814 577898 360986 578134
rect 361222 577898 361394 578134
rect 360814 542454 361394 577898
rect 360814 542218 360986 542454
rect 361222 542218 361394 542454
rect 360814 542134 361394 542218
rect 360814 541898 360986 542134
rect 361222 541898 361394 542134
rect 360814 506454 361394 541898
rect 360814 506218 360986 506454
rect 361222 506218 361394 506454
rect 360814 506134 361394 506218
rect 360814 505898 360986 506134
rect 361222 505898 361394 506134
rect 360814 470454 361394 505898
rect 360814 470218 360986 470454
rect 361222 470218 361394 470454
rect 360814 470134 361394 470218
rect 360814 469898 360986 470134
rect 361222 469898 361394 470134
rect 360814 434454 361394 469898
rect 360814 434218 360986 434454
rect 361222 434218 361394 434454
rect 360814 434134 361394 434218
rect 360814 433898 360986 434134
rect 361222 433898 361394 434134
rect 360814 398454 361394 433898
rect 360814 398218 360986 398454
rect 361222 398218 361394 398454
rect 360814 398134 361394 398218
rect 360814 397898 360986 398134
rect 361222 397898 361394 398134
rect 359595 362948 359661 362949
rect 359595 362884 359596 362948
rect 359660 362884 359661 362948
rect 359595 362883 359661 362884
rect 359598 360858 359658 362883
rect 360814 362454 361394 397898
rect 360814 362218 360986 362454
rect 361222 362218 361394 362454
rect 360814 362134 361394 362218
rect 360814 361898 360986 362134
rect 361222 361898 361394 362134
rect 353254 354658 353426 354894
rect 353662 354658 353834 354894
rect 353254 354574 353834 354658
rect 353254 354338 353426 354574
rect 353662 354338 353834 354574
rect 353254 318894 353834 354338
rect 353254 318658 353426 318894
rect 353662 318658 353834 318894
rect 353254 318574 353834 318658
rect 353254 318338 353426 318574
rect 353662 318338 353834 318574
rect 353254 282894 353834 318338
rect 353254 282658 353426 282894
rect 353662 282658 353834 282894
rect 353254 282574 353834 282658
rect 353254 282338 353426 282574
rect 353662 282338 353834 282574
rect 353254 246894 353834 282338
rect 353254 246658 353426 246894
rect 353662 246658 353834 246894
rect 353254 246574 353834 246658
rect 353254 246338 353426 246574
rect 353662 246338 353834 246574
rect 353254 210894 353834 246338
rect 353254 210658 353426 210894
rect 353662 210658 353834 210894
rect 353254 210574 353834 210658
rect 353254 210338 353426 210574
rect 353662 210338 353834 210574
rect 353254 174894 353834 210338
rect 353254 174658 353426 174894
rect 353662 174658 353834 174894
rect 353254 174574 353834 174658
rect 353254 174338 353426 174574
rect 353662 174338 353834 174574
rect 353254 138894 353834 174338
rect 353254 138658 353426 138894
rect 353662 138658 353834 138894
rect 353254 138574 353834 138658
rect 353254 138338 353426 138574
rect 353662 138338 353834 138574
rect 353254 102894 353834 138338
rect 353254 102658 353426 102894
rect 353662 102658 353834 102894
rect 353254 102574 353834 102658
rect 353254 102338 353426 102574
rect 353662 102338 353834 102574
rect 353254 66894 353834 102338
rect 353254 66658 353426 66894
rect 353662 66658 353834 66894
rect 353254 66574 353834 66658
rect 353254 66338 353426 66574
rect 353662 66338 353834 66574
rect 353254 30894 353834 66338
rect 353254 30658 353426 30894
rect 353662 30658 353834 30894
rect 353254 30574 353834 30658
rect 353254 30338 353426 30574
rect 353662 30338 353834 30574
rect 335254 -6102 335426 -5866
rect 335662 -6102 335834 -5866
rect 335254 -6186 335834 -6102
rect 335254 -6422 335426 -6186
rect 335662 -6422 335834 -6186
rect 335254 -7354 335834 -6422
rect 353254 -6786 353834 30338
rect 360814 326454 361394 361898
rect 360814 326218 360986 326454
rect 361222 326218 361394 326454
rect 360814 326134 361394 326218
rect 360814 325898 360986 326134
rect 361222 325898 361394 326134
rect 360814 290454 361394 325898
rect 360814 290218 360986 290454
rect 361222 290218 361394 290454
rect 360814 290134 361394 290218
rect 360814 289898 360986 290134
rect 361222 289898 361394 290134
rect 360814 254454 361394 289898
rect 360814 254218 360986 254454
rect 361222 254218 361394 254454
rect 360814 254134 361394 254218
rect 360814 253898 360986 254134
rect 361222 253898 361394 254134
rect 360814 218454 361394 253898
rect 360814 218218 360986 218454
rect 361222 218218 361394 218454
rect 360814 218134 361394 218218
rect 360814 217898 360986 218134
rect 361222 217898 361394 218134
rect 360814 182454 361394 217898
rect 360814 182218 360986 182454
rect 361222 182218 361394 182454
rect 360814 182134 361394 182218
rect 360814 181898 360986 182134
rect 361222 181898 361394 182134
rect 360814 146454 361394 181898
rect 360814 146218 360986 146454
rect 361222 146218 361394 146454
rect 360814 146134 361394 146218
rect 360814 145898 360986 146134
rect 361222 145898 361394 146134
rect 360814 110454 361394 145898
rect 360814 110218 360986 110454
rect 361222 110218 361394 110454
rect 360814 110134 361394 110218
rect 360814 109898 360986 110134
rect 361222 109898 361394 110134
rect 360814 74454 361394 109898
rect 360814 74218 360986 74454
rect 361222 74218 361394 74454
rect 360814 74134 361394 74218
rect 360814 73898 360986 74134
rect 361222 73898 361394 74134
rect 360814 38454 361394 73898
rect 360814 38218 360986 38454
rect 361222 38218 361394 38454
rect 360814 38134 361394 38218
rect 360814 37898 360986 38134
rect 361222 37898 361394 38134
rect 360814 2454 361394 37898
rect 360814 2218 360986 2454
rect 361222 2218 361394 2454
rect 360814 2134 361394 2218
rect 360814 1898 360986 2134
rect 361222 1898 361394 2134
rect 360814 -346 361394 1898
rect 360814 -582 360986 -346
rect 361222 -582 361394 -346
rect 360814 -666 361394 -582
rect 360814 -902 360986 -666
rect 361222 -902 361394 -666
rect 360814 -1834 361394 -902
rect 364294 689934 364874 706122
rect 364294 689698 364466 689934
rect 364702 689698 364874 689934
rect 364294 689614 364874 689698
rect 364294 689378 364466 689614
rect 364702 689378 364874 689614
rect 364294 653934 364874 689378
rect 364294 653698 364466 653934
rect 364702 653698 364874 653934
rect 364294 653614 364874 653698
rect 364294 653378 364466 653614
rect 364702 653378 364874 653614
rect 364294 617934 364874 653378
rect 364294 617698 364466 617934
rect 364702 617698 364874 617934
rect 364294 617614 364874 617698
rect 364294 617378 364466 617614
rect 364702 617378 364874 617614
rect 364294 581934 364874 617378
rect 364294 581698 364466 581934
rect 364702 581698 364874 581934
rect 364294 581614 364874 581698
rect 364294 581378 364466 581614
rect 364702 581378 364874 581614
rect 364294 545934 364874 581378
rect 364294 545698 364466 545934
rect 364702 545698 364874 545934
rect 364294 545614 364874 545698
rect 364294 545378 364466 545614
rect 364702 545378 364874 545614
rect 364294 509934 364874 545378
rect 364294 509698 364466 509934
rect 364702 509698 364874 509934
rect 364294 509614 364874 509698
rect 364294 509378 364466 509614
rect 364702 509378 364874 509614
rect 364294 473934 364874 509378
rect 364294 473698 364466 473934
rect 364702 473698 364874 473934
rect 364294 473614 364874 473698
rect 364294 473378 364466 473614
rect 364702 473378 364874 473614
rect 364294 437934 364874 473378
rect 364294 437698 364466 437934
rect 364702 437698 364874 437934
rect 364294 437614 364874 437698
rect 364294 437378 364466 437614
rect 364702 437378 364874 437614
rect 364294 401934 364874 437378
rect 364294 401698 364466 401934
rect 364702 401698 364874 401934
rect 364294 401614 364874 401698
rect 364294 401378 364466 401614
rect 364702 401378 364874 401614
rect 364294 365934 364874 401378
rect 364294 365698 364466 365934
rect 364702 365698 364874 365934
rect 364294 365614 364874 365698
rect 364294 365378 364466 365614
rect 364702 365378 364874 365614
rect 364294 329934 364874 365378
rect 364294 329698 364466 329934
rect 364702 329698 364874 329934
rect 364294 329614 364874 329698
rect 364294 329378 364466 329614
rect 364702 329378 364874 329614
rect 364294 293934 364874 329378
rect 364294 293698 364466 293934
rect 364702 293698 364874 293934
rect 364294 293614 364874 293698
rect 364294 293378 364466 293614
rect 364702 293378 364874 293614
rect 364294 257934 364874 293378
rect 364294 257698 364466 257934
rect 364702 257698 364874 257934
rect 364294 257614 364874 257698
rect 364294 257378 364466 257614
rect 364702 257378 364874 257614
rect 364294 221934 364874 257378
rect 364294 221698 364466 221934
rect 364702 221698 364874 221934
rect 364294 221614 364874 221698
rect 364294 221378 364466 221614
rect 364702 221378 364874 221614
rect 364294 185934 364874 221378
rect 364294 185698 364466 185934
rect 364702 185698 364874 185934
rect 364294 185614 364874 185698
rect 364294 185378 364466 185614
rect 364702 185378 364874 185614
rect 364294 149934 364874 185378
rect 364294 149698 364466 149934
rect 364702 149698 364874 149934
rect 364294 149614 364874 149698
rect 364294 149378 364466 149614
rect 364702 149378 364874 149614
rect 364294 113934 364874 149378
rect 364294 113698 364466 113934
rect 364702 113698 364874 113934
rect 364294 113614 364874 113698
rect 364294 113378 364466 113614
rect 364702 113378 364874 113614
rect 364294 77934 364874 113378
rect 364294 77698 364466 77934
rect 364702 77698 364874 77934
rect 364294 77614 364874 77698
rect 364294 77378 364466 77614
rect 364702 77378 364874 77614
rect 364294 41934 364874 77378
rect 364294 41698 364466 41934
rect 364702 41698 364874 41934
rect 364294 41614 364874 41698
rect 364294 41378 364466 41614
rect 364702 41378 364874 41614
rect 364294 5934 364874 41378
rect 364294 5698 364466 5934
rect 364702 5698 364874 5934
rect 364294 5614 364874 5698
rect 364294 5378 364466 5614
rect 364702 5378 364874 5614
rect 364294 -2186 364874 5378
rect 364294 -2422 364466 -2186
rect 364702 -2422 364874 -2186
rect 364294 -2506 364874 -2422
rect 364294 -2742 364466 -2506
rect 364702 -2742 364874 -2506
rect 364294 -3674 364874 -2742
rect 367774 693414 368354 707962
rect 367774 693178 367946 693414
rect 368182 693178 368354 693414
rect 367774 693094 368354 693178
rect 367774 692858 367946 693094
rect 368182 692858 368354 693094
rect 367774 657414 368354 692858
rect 367774 657178 367946 657414
rect 368182 657178 368354 657414
rect 367774 657094 368354 657178
rect 367774 656858 367946 657094
rect 368182 656858 368354 657094
rect 367774 621414 368354 656858
rect 367774 621178 367946 621414
rect 368182 621178 368354 621414
rect 367774 621094 368354 621178
rect 367774 620858 367946 621094
rect 368182 620858 368354 621094
rect 367774 585414 368354 620858
rect 367774 585178 367946 585414
rect 368182 585178 368354 585414
rect 367774 585094 368354 585178
rect 367774 584858 367946 585094
rect 368182 584858 368354 585094
rect 367774 549414 368354 584858
rect 367774 549178 367946 549414
rect 368182 549178 368354 549414
rect 367774 549094 368354 549178
rect 367774 548858 367946 549094
rect 368182 548858 368354 549094
rect 367774 513414 368354 548858
rect 367774 513178 367946 513414
rect 368182 513178 368354 513414
rect 367774 513094 368354 513178
rect 367774 512858 367946 513094
rect 368182 512858 368354 513094
rect 367774 477414 368354 512858
rect 367774 477178 367946 477414
rect 368182 477178 368354 477414
rect 367774 477094 368354 477178
rect 367774 476858 367946 477094
rect 368182 476858 368354 477094
rect 367774 441414 368354 476858
rect 367774 441178 367946 441414
rect 368182 441178 368354 441414
rect 367774 441094 368354 441178
rect 367774 440858 367946 441094
rect 368182 440858 368354 441094
rect 367774 405414 368354 440858
rect 367774 405178 367946 405414
rect 368182 405178 368354 405414
rect 367774 405094 368354 405178
rect 367774 404858 367946 405094
rect 368182 404858 368354 405094
rect 367774 369414 368354 404858
rect 367774 369178 367946 369414
rect 368182 369178 368354 369414
rect 367774 369094 368354 369178
rect 367774 368858 367946 369094
rect 368182 368858 368354 369094
rect 367774 333414 368354 368858
rect 367774 333178 367946 333414
rect 368182 333178 368354 333414
rect 367774 333094 368354 333178
rect 367774 332858 367946 333094
rect 368182 332858 368354 333094
rect 367774 297414 368354 332858
rect 367774 297178 367946 297414
rect 368182 297178 368354 297414
rect 367774 297094 368354 297178
rect 367774 296858 367946 297094
rect 368182 296858 368354 297094
rect 367774 261414 368354 296858
rect 367774 261178 367946 261414
rect 368182 261178 368354 261414
rect 367774 261094 368354 261178
rect 367774 260858 367946 261094
rect 368182 260858 368354 261094
rect 367774 225414 368354 260858
rect 367774 225178 367946 225414
rect 368182 225178 368354 225414
rect 367774 225094 368354 225178
rect 367774 224858 367946 225094
rect 368182 224858 368354 225094
rect 367774 189414 368354 224858
rect 367774 189178 367946 189414
rect 368182 189178 368354 189414
rect 367774 189094 368354 189178
rect 367774 188858 367946 189094
rect 368182 188858 368354 189094
rect 367774 153414 368354 188858
rect 367774 153178 367946 153414
rect 368182 153178 368354 153414
rect 367774 153094 368354 153178
rect 367774 152858 367946 153094
rect 368182 152858 368354 153094
rect 367774 117414 368354 152858
rect 367774 117178 367946 117414
rect 368182 117178 368354 117414
rect 367774 117094 368354 117178
rect 367774 116858 367946 117094
rect 368182 116858 368354 117094
rect 367774 81414 368354 116858
rect 367774 81178 367946 81414
rect 368182 81178 368354 81414
rect 367774 81094 368354 81178
rect 367774 80858 367946 81094
rect 368182 80858 368354 81094
rect 367774 45414 368354 80858
rect 367774 45178 367946 45414
rect 368182 45178 368354 45414
rect 367774 45094 368354 45178
rect 367774 44858 367946 45094
rect 368182 44858 368354 45094
rect 367774 9414 368354 44858
rect 367774 9178 367946 9414
rect 368182 9178 368354 9414
rect 367774 9094 368354 9178
rect 367774 8858 367946 9094
rect 368182 8858 368354 9094
rect 367774 -4026 368354 8858
rect 367774 -4262 367946 -4026
rect 368182 -4262 368354 -4026
rect 367774 -4346 368354 -4262
rect 367774 -4582 367946 -4346
rect 368182 -4582 368354 -4346
rect 367774 -5514 368354 -4582
rect 371254 696894 371834 709802
rect 389254 711278 389834 711290
rect 389254 711042 389426 711278
rect 389662 711042 389834 711278
rect 389254 710958 389834 711042
rect 389254 710722 389426 710958
rect 389662 710722 389834 710958
rect 385774 709438 386354 709450
rect 385774 709202 385946 709438
rect 386182 709202 386354 709438
rect 385774 709118 386354 709202
rect 385774 708882 385946 709118
rect 386182 708882 386354 709118
rect 382294 707598 382874 707610
rect 382294 707362 382466 707598
rect 382702 707362 382874 707598
rect 382294 707278 382874 707362
rect 382294 707042 382466 707278
rect 382702 707042 382874 707278
rect 371254 696658 371426 696894
rect 371662 696658 371834 696894
rect 371254 696574 371834 696658
rect 371254 696338 371426 696574
rect 371662 696338 371834 696574
rect 371254 660894 371834 696338
rect 371254 660658 371426 660894
rect 371662 660658 371834 660894
rect 371254 660574 371834 660658
rect 371254 660338 371426 660574
rect 371662 660338 371834 660574
rect 371254 624894 371834 660338
rect 371254 624658 371426 624894
rect 371662 624658 371834 624894
rect 371254 624574 371834 624658
rect 371254 624338 371426 624574
rect 371662 624338 371834 624574
rect 371254 588894 371834 624338
rect 371254 588658 371426 588894
rect 371662 588658 371834 588894
rect 371254 588574 371834 588658
rect 371254 588338 371426 588574
rect 371662 588338 371834 588574
rect 371254 552894 371834 588338
rect 371254 552658 371426 552894
rect 371662 552658 371834 552894
rect 371254 552574 371834 552658
rect 371254 552338 371426 552574
rect 371662 552338 371834 552574
rect 371254 516894 371834 552338
rect 371254 516658 371426 516894
rect 371662 516658 371834 516894
rect 371254 516574 371834 516658
rect 371254 516338 371426 516574
rect 371662 516338 371834 516574
rect 371254 480894 371834 516338
rect 371254 480658 371426 480894
rect 371662 480658 371834 480894
rect 371254 480574 371834 480658
rect 371254 480338 371426 480574
rect 371662 480338 371834 480574
rect 371254 444894 371834 480338
rect 371254 444658 371426 444894
rect 371662 444658 371834 444894
rect 371254 444574 371834 444658
rect 371254 444338 371426 444574
rect 371662 444338 371834 444574
rect 371254 408894 371834 444338
rect 371254 408658 371426 408894
rect 371662 408658 371834 408894
rect 371254 408574 371834 408658
rect 371254 408338 371426 408574
rect 371662 408338 371834 408574
rect 371254 372894 371834 408338
rect 371254 372658 371426 372894
rect 371662 372658 371834 372894
rect 371254 372574 371834 372658
rect 371254 372338 371426 372574
rect 371662 372338 371834 372574
rect 371254 336894 371834 372338
rect 371254 336658 371426 336894
rect 371662 336658 371834 336894
rect 371254 336574 371834 336658
rect 371254 336338 371426 336574
rect 371662 336338 371834 336574
rect 371254 300894 371834 336338
rect 371254 300658 371426 300894
rect 371662 300658 371834 300894
rect 371254 300574 371834 300658
rect 371254 300338 371426 300574
rect 371662 300338 371834 300574
rect 371254 264894 371834 300338
rect 371254 264658 371426 264894
rect 371662 264658 371834 264894
rect 371254 264574 371834 264658
rect 371254 264338 371426 264574
rect 371662 264338 371834 264574
rect 371254 228894 371834 264338
rect 371254 228658 371426 228894
rect 371662 228658 371834 228894
rect 371254 228574 371834 228658
rect 371254 228338 371426 228574
rect 371662 228338 371834 228574
rect 371254 192894 371834 228338
rect 371254 192658 371426 192894
rect 371662 192658 371834 192894
rect 371254 192574 371834 192658
rect 371254 192338 371426 192574
rect 371662 192338 371834 192574
rect 371254 156894 371834 192338
rect 371254 156658 371426 156894
rect 371662 156658 371834 156894
rect 371254 156574 371834 156658
rect 371254 156338 371426 156574
rect 371662 156338 371834 156574
rect 371254 120894 371834 156338
rect 371254 120658 371426 120894
rect 371662 120658 371834 120894
rect 371254 120574 371834 120658
rect 371254 120338 371426 120574
rect 371662 120338 371834 120574
rect 371254 84894 371834 120338
rect 371254 84658 371426 84894
rect 371662 84658 371834 84894
rect 371254 84574 371834 84658
rect 371254 84338 371426 84574
rect 371662 84338 371834 84574
rect 371254 48894 371834 84338
rect 371254 48658 371426 48894
rect 371662 48658 371834 48894
rect 371254 48574 371834 48658
rect 371254 48338 371426 48574
rect 371662 48338 371834 48574
rect 371254 12894 371834 48338
rect 371254 12658 371426 12894
rect 371662 12658 371834 12894
rect 371254 12574 371834 12658
rect 371254 12338 371426 12574
rect 371662 12338 371834 12574
rect 353254 -7022 353426 -6786
rect 353662 -7022 353834 -6786
rect 353254 -7106 353834 -7022
rect 353254 -7342 353426 -7106
rect 353662 -7342 353834 -7106
rect 353254 -7354 353834 -7342
rect 371254 -5866 371834 12338
rect 378814 705758 379394 705770
rect 378814 705522 378986 705758
rect 379222 705522 379394 705758
rect 378814 705438 379394 705522
rect 378814 705202 378986 705438
rect 379222 705202 379394 705438
rect 378814 668454 379394 705202
rect 378814 668218 378986 668454
rect 379222 668218 379394 668454
rect 378814 668134 379394 668218
rect 378814 667898 378986 668134
rect 379222 667898 379394 668134
rect 378814 632454 379394 667898
rect 378814 632218 378986 632454
rect 379222 632218 379394 632454
rect 378814 632134 379394 632218
rect 378814 631898 378986 632134
rect 379222 631898 379394 632134
rect 378814 596454 379394 631898
rect 378814 596218 378986 596454
rect 379222 596218 379394 596454
rect 378814 596134 379394 596218
rect 378814 595898 378986 596134
rect 379222 595898 379394 596134
rect 378814 560454 379394 595898
rect 378814 560218 378986 560454
rect 379222 560218 379394 560454
rect 378814 560134 379394 560218
rect 378814 559898 378986 560134
rect 379222 559898 379394 560134
rect 378814 524454 379394 559898
rect 378814 524218 378986 524454
rect 379222 524218 379394 524454
rect 378814 524134 379394 524218
rect 378814 523898 378986 524134
rect 379222 523898 379394 524134
rect 378814 488454 379394 523898
rect 378814 488218 378986 488454
rect 379222 488218 379394 488454
rect 378814 488134 379394 488218
rect 378814 487898 378986 488134
rect 379222 487898 379394 488134
rect 378814 452454 379394 487898
rect 378814 452218 378986 452454
rect 379222 452218 379394 452454
rect 378814 452134 379394 452218
rect 378814 451898 378986 452134
rect 379222 451898 379394 452134
rect 378814 416454 379394 451898
rect 378814 416218 378986 416454
rect 379222 416218 379394 416454
rect 378814 416134 379394 416218
rect 378814 415898 378986 416134
rect 379222 415898 379394 416134
rect 378814 380454 379394 415898
rect 378814 380218 378986 380454
rect 379222 380218 379394 380454
rect 378814 380134 379394 380218
rect 378814 379898 378986 380134
rect 379222 379898 379394 380134
rect 378814 344454 379394 379898
rect 378814 344218 378986 344454
rect 379222 344218 379394 344454
rect 378814 344134 379394 344218
rect 378814 343898 378986 344134
rect 379222 343898 379394 344134
rect 378814 308454 379394 343898
rect 378814 308218 378986 308454
rect 379222 308218 379394 308454
rect 378814 308134 379394 308218
rect 378814 307898 378986 308134
rect 379222 307898 379394 308134
rect 378814 272454 379394 307898
rect 378814 272218 378986 272454
rect 379222 272218 379394 272454
rect 378814 272134 379394 272218
rect 378814 271898 378986 272134
rect 379222 271898 379394 272134
rect 378814 236454 379394 271898
rect 378814 236218 378986 236454
rect 379222 236218 379394 236454
rect 378814 236134 379394 236218
rect 378814 235898 378986 236134
rect 379222 235898 379394 236134
rect 378814 200454 379394 235898
rect 378814 200218 378986 200454
rect 379222 200218 379394 200454
rect 378814 200134 379394 200218
rect 378814 199898 378986 200134
rect 379222 199898 379394 200134
rect 378814 164454 379394 199898
rect 378814 164218 378986 164454
rect 379222 164218 379394 164454
rect 378814 164134 379394 164218
rect 378814 163898 378986 164134
rect 379222 163898 379394 164134
rect 378814 128454 379394 163898
rect 378814 128218 378986 128454
rect 379222 128218 379394 128454
rect 378814 128134 379394 128218
rect 378814 127898 378986 128134
rect 379222 127898 379394 128134
rect 378814 92454 379394 127898
rect 378814 92218 378986 92454
rect 379222 92218 379394 92454
rect 378814 92134 379394 92218
rect 378814 91898 378986 92134
rect 379222 91898 379394 92134
rect 378814 56454 379394 91898
rect 378814 56218 378986 56454
rect 379222 56218 379394 56454
rect 378814 56134 379394 56218
rect 378814 55898 378986 56134
rect 379222 55898 379394 56134
rect 378814 20454 379394 55898
rect 378814 20218 378986 20454
rect 379222 20218 379394 20454
rect 378814 20134 379394 20218
rect 378814 19898 378986 20134
rect 379222 19898 379394 20134
rect 378814 -1266 379394 19898
rect 378814 -1502 378986 -1266
rect 379222 -1502 379394 -1266
rect 378814 -1586 379394 -1502
rect 378814 -1822 378986 -1586
rect 379222 -1822 379394 -1586
rect 378814 -1834 379394 -1822
rect 382294 671934 382874 707042
rect 382294 671698 382466 671934
rect 382702 671698 382874 671934
rect 382294 671614 382874 671698
rect 382294 671378 382466 671614
rect 382702 671378 382874 671614
rect 382294 635934 382874 671378
rect 382294 635698 382466 635934
rect 382702 635698 382874 635934
rect 382294 635614 382874 635698
rect 382294 635378 382466 635614
rect 382702 635378 382874 635614
rect 382294 599934 382874 635378
rect 382294 599698 382466 599934
rect 382702 599698 382874 599934
rect 382294 599614 382874 599698
rect 382294 599378 382466 599614
rect 382702 599378 382874 599614
rect 382294 563934 382874 599378
rect 382294 563698 382466 563934
rect 382702 563698 382874 563934
rect 382294 563614 382874 563698
rect 382294 563378 382466 563614
rect 382702 563378 382874 563614
rect 382294 527934 382874 563378
rect 382294 527698 382466 527934
rect 382702 527698 382874 527934
rect 382294 527614 382874 527698
rect 382294 527378 382466 527614
rect 382702 527378 382874 527614
rect 382294 491934 382874 527378
rect 382294 491698 382466 491934
rect 382702 491698 382874 491934
rect 382294 491614 382874 491698
rect 382294 491378 382466 491614
rect 382702 491378 382874 491614
rect 382294 455934 382874 491378
rect 382294 455698 382466 455934
rect 382702 455698 382874 455934
rect 382294 455614 382874 455698
rect 382294 455378 382466 455614
rect 382702 455378 382874 455614
rect 382294 419934 382874 455378
rect 382294 419698 382466 419934
rect 382702 419698 382874 419934
rect 382294 419614 382874 419698
rect 382294 419378 382466 419614
rect 382702 419378 382874 419614
rect 382294 383934 382874 419378
rect 382294 383698 382466 383934
rect 382702 383698 382874 383934
rect 382294 383614 382874 383698
rect 382294 383378 382466 383614
rect 382702 383378 382874 383614
rect 382294 347934 382874 383378
rect 382294 347698 382466 347934
rect 382702 347698 382874 347934
rect 382294 347614 382874 347698
rect 382294 347378 382466 347614
rect 382702 347378 382874 347614
rect 382294 311934 382874 347378
rect 382294 311698 382466 311934
rect 382702 311698 382874 311934
rect 382294 311614 382874 311698
rect 382294 311378 382466 311614
rect 382702 311378 382874 311614
rect 382294 275934 382874 311378
rect 382294 275698 382466 275934
rect 382702 275698 382874 275934
rect 382294 275614 382874 275698
rect 382294 275378 382466 275614
rect 382702 275378 382874 275614
rect 382294 239934 382874 275378
rect 382294 239698 382466 239934
rect 382702 239698 382874 239934
rect 382294 239614 382874 239698
rect 382294 239378 382466 239614
rect 382702 239378 382874 239614
rect 382294 203934 382874 239378
rect 382294 203698 382466 203934
rect 382702 203698 382874 203934
rect 382294 203614 382874 203698
rect 382294 203378 382466 203614
rect 382702 203378 382874 203614
rect 382294 167934 382874 203378
rect 382294 167698 382466 167934
rect 382702 167698 382874 167934
rect 382294 167614 382874 167698
rect 382294 167378 382466 167614
rect 382702 167378 382874 167614
rect 382294 131934 382874 167378
rect 382294 131698 382466 131934
rect 382702 131698 382874 131934
rect 382294 131614 382874 131698
rect 382294 131378 382466 131614
rect 382702 131378 382874 131614
rect 382294 95934 382874 131378
rect 382294 95698 382466 95934
rect 382702 95698 382874 95934
rect 382294 95614 382874 95698
rect 382294 95378 382466 95614
rect 382702 95378 382874 95614
rect 382294 59934 382874 95378
rect 382294 59698 382466 59934
rect 382702 59698 382874 59934
rect 382294 59614 382874 59698
rect 382294 59378 382466 59614
rect 382702 59378 382874 59614
rect 382294 23934 382874 59378
rect 382294 23698 382466 23934
rect 382702 23698 382874 23934
rect 382294 23614 382874 23698
rect 382294 23378 382466 23614
rect 382702 23378 382874 23614
rect 382294 -3106 382874 23378
rect 382294 -3342 382466 -3106
rect 382702 -3342 382874 -3106
rect 382294 -3426 382874 -3342
rect 382294 -3662 382466 -3426
rect 382702 -3662 382874 -3426
rect 382294 -3674 382874 -3662
rect 385774 675414 386354 708882
rect 385774 675178 385946 675414
rect 386182 675178 386354 675414
rect 385774 675094 386354 675178
rect 385774 674858 385946 675094
rect 386182 674858 386354 675094
rect 385774 639414 386354 674858
rect 385774 639178 385946 639414
rect 386182 639178 386354 639414
rect 385774 639094 386354 639178
rect 385774 638858 385946 639094
rect 386182 638858 386354 639094
rect 385774 603414 386354 638858
rect 385774 603178 385946 603414
rect 386182 603178 386354 603414
rect 385774 603094 386354 603178
rect 385774 602858 385946 603094
rect 386182 602858 386354 603094
rect 385774 567414 386354 602858
rect 385774 567178 385946 567414
rect 386182 567178 386354 567414
rect 385774 567094 386354 567178
rect 385774 566858 385946 567094
rect 386182 566858 386354 567094
rect 385774 531414 386354 566858
rect 385774 531178 385946 531414
rect 386182 531178 386354 531414
rect 385774 531094 386354 531178
rect 385774 530858 385946 531094
rect 386182 530858 386354 531094
rect 385774 495414 386354 530858
rect 385774 495178 385946 495414
rect 386182 495178 386354 495414
rect 385774 495094 386354 495178
rect 385774 494858 385946 495094
rect 386182 494858 386354 495094
rect 385774 459414 386354 494858
rect 385774 459178 385946 459414
rect 386182 459178 386354 459414
rect 385774 459094 386354 459178
rect 385774 458858 385946 459094
rect 386182 458858 386354 459094
rect 385774 423414 386354 458858
rect 385774 423178 385946 423414
rect 386182 423178 386354 423414
rect 385774 423094 386354 423178
rect 385774 422858 385946 423094
rect 386182 422858 386354 423094
rect 385774 387414 386354 422858
rect 385774 387178 385946 387414
rect 386182 387178 386354 387414
rect 385774 387094 386354 387178
rect 385774 386858 385946 387094
rect 386182 386858 386354 387094
rect 385774 351414 386354 386858
rect 385774 351178 385946 351414
rect 386182 351178 386354 351414
rect 385774 351094 386354 351178
rect 385774 350858 385946 351094
rect 386182 350858 386354 351094
rect 385774 315414 386354 350858
rect 385774 315178 385946 315414
rect 386182 315178 386354 315414
rect 385774 315094 386354 315178
rect 385774 314858 385946 315094
rect 386182 314858 386354 315094
rect 385774 279414 386354 314858
rect 385774 279178 385946 279414
rect 386182 279178 386354 279414
rect 385774 279094 386354 279178
rect 385774 278858 385946 279094
rect 386182 278858 386354 279094
rect 385774 243414 386354 278858
rect 385774 243178 385946 243414
rect 386182 243178 386354 243414
rect 385774 243094 386354 243178
rect 385774 242858 385946 243094
rect 386182 242858 386354 243094
rect 385774 207414 386354 242858
rect 385774 207178 385946 207414
rect 386182 207178 386354 207414
rect 385774 207094 386354 207178
rect 385774 206858 385946 207094
rect 386182 206858 386354 207094
rect 385774 171414 386354 206858
rect 385774 171178 385946 171414
rect 386182 171178 386354 171414
rect 385774 171094 386354 171178
rect 385774 170858 385946 171094
rect 386182 170858 386354 171094
rect 385774 135414 386354 170858
rect 385774 135178 385946 135414
rect 386182 135178 386354 135414
rect 385774 135094 386354 135178
rect 385774 134858 385946 135094
rect 386182 134858 386354 135094
rect 385774 99414 386354 134858
rect 385774 99178 385946 99414
rect 386182 99178 386354 99414
rect 385774 99094 386354 99178
rect 385774 98858 385946 99094
rect 386182 98858 386354 99094
rect 385774 63414 386354 98858
rect 385774 63178 385946 63414
rect 386182 63178 386354 63414
rect 385774 63094 386354 63178
rect 385774 62858 385946 63094
rect 386182 62858 386354 63094
rect 385774 27414 386354 62858
rect 385774 27178 385946 27414
rect 386182 27178 386354 27414
rect 385774 27094 386354 27178
rect 385774 26858 385946 27094
rect 386182 26858 386354 27094
rect 385774 -4946 386354 26858
rect 385774 -5182 385946 -4946
rect 386182 -5182 386354 -4946
rect 385774 -5266 386354 -5182
rect 385774 -5502 385946 -5266
rect 386182 -5502 386354 -5266
rect 385774 -5514 386354 -5502
rect 389254 678894 389834 710722
rect 407254 710358 407834 711290
rect 407254 710122 407426 710358
rect 407662 710122 407834 710358
rect 407254 710038 407834 710122
rect 407254 709802 407426 710038
rect 407662 709802 407834 710038
rect 403774 708518 404354 709450
rect 403774 708282 403946 708518
rect 404182 708282 404354 708518
rect 403774 708198 404354 708282
rect 403774 707962 403946 708198
rect 404182 707962 404354 708198
rect 400294 706678 400874 707610
rect 400294 706442 400466 706678
rect 400702 706442 400874 706678
rect 400294 706358 400874 706442
rect 400294 706122 400466 706358
rect 400702 706122 400874 706358
rect 389254 678658 389426 678894
rect 389662 678658 389834 678894
rect 389254 678574 389834 678658
rect 389254 678338 389426 678574
rect 389662 678338 389834 678574
rect 389254 642894 389834 678338
rect 389254 642658 389426 642894
rect 389662 642658 389834 642894
rect 389254 642574 389834 642658
rect 389254 642338 389426 642574
rect 389662 642338 389834 642574
rect 389254 606894 389834 642338
rect 389254 606658 389426 606894
rect 389662 606658 389834 606894
rect 389254 606574 389834 606658
rect 389254 606338 389426 606574
rect 389662 606338 389834 606574
rect 389254 570894 389834 606338
rect 389254 570658 389426 570894
rect 389662 570658 389834 570894
rect 389254 570574 389834 570658
rect 389254 570338 389426 570574
rect 389662 570338 389834 570574
rect 389254 534894 389834 570338
rect 389254 534658 389426 534894
rect 389662 534658 389834 534894
rect 389254 534574 389834 534658
rect 389254 534338 389426 534574
rect 389662 534338 389834 534574
rect 389254 498894 389834 534338
rect 389254 498658 389426 498894
rect 389662 498658 389834 498894
rect 389254 498574 389834 498658
rect 389254 498338 389426 498574
rect 389662 498338 389834 498574
rect 389254 462894 389834 498338
rect 389254 462658 389426 462894
rect 389662 462658 389834 462894
rect 389254 462574 389834 462658
rect 389254 462338 389426 462574
rect 389662 462338 389834 462574
rect 389254 426894 389834 462338
rect 389254 426658 389426 426894
rect 389662 426658 389834 426894
rect 389254 426574 389834 426658
rect 389254 426338 389426 426574
rect 389662 426338 389834 426574
rect 389254 390894 389834 426338
rect 389254 390658 389426 390894
rect 389662 390658 389834 390894
rect 389254 390574 389834 390658
rect 389254 390338 389426 390574
rect 389662 390338 389834 390574
rect 389254 354894 389834 390338
rect 389254 354658 389426 354894
rect 389662 354658 389834 354894
rect 389254 354574 389834 354658
rect 389254 354338 389426 354574
rect 389662 354338 389834 354574
rect 389254 318894 389834 354338
rect 389254 318658 389426 318894
rect 389662 318658 389834 318894
rect 389254 318574 389834 318658
rect 389254 318338 389426 318574
rect 389662 318338 389834 318574
rect 389254 282894 389834 318338
rect 389254 282658 389426 282894
rect 389662 282658 389834 282894
rect 389254 282574 389834 282658
rect 389254 282338 389426 282574
rect 389662 282338 389834 282574
rect 389254 246894 389834 282338
rect 389254 246658 389426 246894
rect 389662 246658 389834 246894
rect 389254 246574 389834 246658
rect 389254 246338 389426 246574
rect 389662 246338 389834 246574
rect 389254 210894 389834 246338
rect 389254 210658 389426 210894
rect 389662 210658 389834 210894
rect 389254 210574 389834 210658
rect 389254 210338 389426 210574
rect 389662 210338 389834 210574
rect 389254 174894 389834 210338
rect 389254 174658 389426 174894
rect 389662 174658 389834 174894
rect 389254 174574 389834 174658
rect 389254 174338 389426 174574
rect 389662 174338 389834 174574
rect 389254 138894 389834 174338
rect 389254 138658 389426 138894
rect 389662 138658 389834 138894
rect 389254 138574 389834 138658
rect 389254 138338 389426 138574
rect 389662 138338 389834 138574
rect 389254 102894 389834 138338
rect 389254 102658 389426 102894
rect 389662 102658 389834 102894
rect 389254 102574 389834 102658
rect 389254 102338 389426 102574
rect 389662 102338 389834 102574
rect 389254 66894 389834 102338
rect 389254 66658 389426 66894
rect 389662 66658 389834 66894
rect 389254 66574 389834 66658
rect 389254 66338 389426 66574
rect 389662 66338 389834 66574
rect 389254 30894 389834 66338
rect 389254 30658 389426 30894
rect 389662 30658 389834 30894
rect 389254 30574 389834 30658
rect 389254 30338 389426 30574
rect 389662 30338 389834 30574
rect 371254 -6102 371426 -5866
rect 371662 -6102 371834 -5866
rect 371254 -6186 371834 -6102
rect 371254 -6422 371426 -6186
rect 371662 -6422 371834 -6186
rect 371254 -7354 371834 -6422
rect 389254 -6786 389834 30338
rect 396814 704838 397394 705770
rect 396814 704602 396986 704838
rect 397222 704602 397394 704838
rect 396814 704518 397394 704602
rect 396814 704282 396986 704518
rect 397222 704282 397394 704518
rect 396814 686454 397394 704282
rect 396814 686218 396986 686454
rect 397222 686218 397394 686454
rect 396814 686134 397394 686218
rect 396814 685898 396986 686134
rect 397222 685898 397394 686134
rect 396814 650454 397394 685898
rect 396814 650218 396986 650454
rect 397222 650218 397394 650454
rect 396814 650134 397394 650218
rect 396814 649898 396986 650134
rect 397222 649898 397394 650134
rect 396814 614454 397394 649898
rect 396814 614218 396986 614454
rect 397222 614218 397394 614454
rect 396814 614134 397394 614218
rect 396814 613898 396986 614134
rect 397222 613898 397394 614134
rect 396814 578454 397394 613898
rect 396814 578218 396986 578454
rect 397222 578218 397394 578454
rect 396814 578134 397394 578218
rect 396814 577898 396986 578134
rect 397222 577898 397394 578134
rect 396814 542454 397394 577898
rect 396814 542218 396986 542454
rect 397222 542218 397394 542454
rect 396814 542134 397394 542218
rect 396814 541898 396986 542134
rect 397222 541898 397394 542134
rect 396814 506454 397394 541898
rect 396814 506218 396986 506454
rect 397222 506218 397394 506454
rect 396814 506134 397394 506218
rect 396814 505898 396986 506134
rect 397222 505898 397394 506134
rect 396814 470454 397394 505898
rect 396814 470218 396986 470454
rect 397222 470218 397394 470454
rect 396814 470134 397394 470218
rect 396814 469898 396986 470134
rect 397222 469898 397394 470134
rect 396814 434454 397394 469898
rect 396814 434218 396986 434454
rect 397222 434218 397394 434454
rect 396814 434134 397394 434218
rect 396814 433898 396986 434134
rect 397222 433898 397394 434134
rect 396814 398454 397394 433898
rect 396814 398218 396986 398454
rect 397222 398218 397394 398454
rect 396814 398134 397394 398218
rect 396814 397898 396986 398134
rect 397222 397898 397394 398134
rect 396814 362454 397394 397898
rect 396814 362218 396986 362454
rect 397222 362218 397394 362454
rect 396814 362134 397394 362218
rect 396814 361898 396986 362134
rect 397222 361898 397394 362134
rect 396814 326454 397394 361898
rect 396814 326218 396986 326454
rect 397222 326218 397394 326454
rect 396814 326134 397394 326218
rect 396814 325898 396986 326134
rect 397222 325898 397394 326134
rect 396814 290454 397394 325898
rect 396814 290218 396986 290454
rect 397222 290218 397394 290454
rect 396814 290134 397394 290218
rect 396814 289898 396986 290134
rect 397222 289898 397394 290134
rect 396814 254454 397394 289898
rect 396814 254218 396986 254454
rect 397222 254218 397394 254454
rect 396814 254134 397394 254218
rect 396814 253898 396986 254134
rect 397222 253898 397394 254134
rect 396814 218454 397394 253898
rect 396814 218218 396986 218454
rect 397222 218218 397394 218454
rect 396814 218134 397394 218218
rect 396814 217898 396986 218134
rect 397222 217898 397394 218134
rect 396814 182454 397394 217898
rect 396814 182218 396986 182454
rect 397222 182218 397394 182454
rect 396814 182134 397394 182218
rect 396814 181898 396986 182134
rect 397222 181898 397394 182134
rect 396814 146454 397394 181898
rect 396814 146218 396986 146454
rect 397222 146218 397394 146454
rect 396814 146134 397394 146218
rect 396814 145898 396986 146134
rect 397222 145898 397394 146134
rect 396814 110454 397394 145898
rect 396814 110218 396986 110454
rect 397222 110218 397394 110454
rect 396814 110134 397394 110218
rect 396814 109898 396986 110134
rect 397222 109898 397394 110134
rect 396814 74454 397394 109898
rect 396814 74218 396986 74454
rect 397222 74218 397394 74454
rect 396814 74134 397394 74218
rect 396814 73898 396986 74134
rect 397222 73898 397394 74134
rect 396814 38454 397394 73898
rect 396814 38218 396986 38454
rect 397222 38218 397394 38454
rect 396814 38134 397394 38218
rect 396814 37898 396986 38134
rect 397222 37898 397394 38134
rect 396814 2454 397394 37898
rect 396814 2218 396986 2454
rect 397222 2218 397394 2454
rect 396814 2134 397394 2218
rect 396814 1898 396986 2134
rect 397222 1898 397394 2134
rect 396814 -346 397394 1898
rect 396814 -582 396986 -346
rect 397222 -582 397394 -346
rect 396814 -666 397394 -582
rect 396814 -902 396986 -666
rect 397222 -902 397394 -666
rect 396814 -1834 397394 -902
rect 400294 689934 400874 706122
rect 400294 689698 400466 689934
rect 400702 689698 400874 689934
rect 400294 689614 400874 689698
rect 400294 689378 400466 689614
rect 400702 689378 400874 689614
rect 400294 653934 400874 689378
rect 400294 653698 400466 653934
rect 400702 653698 400874 653934
rect 400294 653614 400874 653698
rect 400294 653378 400466 653614
rect 400702 653378 400874 653614
rect 400294 617934 400874 653378
rect 400294 617698 400466 617934
rect 400702 617698 400874 617934
rect 400294 617614 400874 617698
rect 400294 617378 400466 617614
rect 400702 617378 400874 617614
rect 400294 581934 400874 617378
rect 400294 581698 400466 581934
rect 400702 581698 400874 581934
rect 400294 581614 400874 581698
rect 400294 581378 400466 581614
rect 400702 581378 400874 581614
rect 400294 545934 400874 581378
rect 400294 545698 400466 545934
rect 400702 545698 400874 545934
rect 400294 545614 400874 545698
rect 400294 545378 400466 545614
rect 400702 545378 400874 545614
rect 400294 509934 400874 545378
rect 400294 509698 400466 509934
rect 400702 509698 400874 509934
rect 400294 509614 400874 509698
rect 400294 509378 400466 509614
rect 400702 509378 400874 509614
rect 400294 473934 400874 509378
rect 400294 473698 400466 473934
rect 400702 473698 400874 473934
rect 400294 473614 400874 473698
rect 400294 473378 400466 473614
rect 400702 473378 400874 473614
rect 400294 437934 400874 473378
rect 400294 437698 400466 437934
rect 400702 437698 400874 437934
rect 400294 437614 400874 437698
rect 400294 437378 400466 437614
rect 400702 437378 400874 437614
rect 400294 401934 400874 437378
rect 400294 401698 400466 401934
rect 400702 401698 400874 401934
rect 400294 401614 400874 401698
rect 400294 401378 400466 401614
rect 400702 401378 400874 401614
rect 400294 365934 400874 401378
rect 400294 365698 400466 365934
rect 400702 365698 400874 365934
rect 400294 365614 400874 365698
rect 400294 365378 400466 365614
rect 400702 365378 400874 365614
rect 400294 329934 400874 365378
rect 400294 329698 400466 329934
rect 400702 329698 400874 329934
rect 400294 329614 400874 329698
rect 400294 329378 400466 329614
rect 400702 329378 400874 329614
rect 400294 293934 400874 329378
rect 400294 293698 400466 293934
rect 400702 293698 400874 293934
rect 400294 293614 400874 293698
rect 400294 293378 400466 293614
rect 400702 293378 400874 293614
rect 400294 257934 400874 293378
rect 400294 257698 400466 257934
rect 400702 257698 400874 257934
rect 400294 257614 400874 257698
rect 400294 257378 400466 257614
rect 400702 257378 400874 257614
rect 400294 221934 400874 257378
rect 400294 221698 400466 221934
rect 400702 221698 400874 221934
rect 400294 221614 400874 221698
rect 400294 221378 400466 221614
rect 400702 221378 400874 221614
rect 400294 185934 400874 221378
rect 400294 185698 400466 185934
rect 400702 185698 400874 185934
rect 400294 185614 400874 185698
rect 400294 185378 400466 185614
rect 400702 185378 400874 185614
rect 400294 149934 400874 185378
rect 400294 149698 400466 149934
rect 400702 149698 400874 149934
rect 400294 149614 400874 149698
rect 400294 149378 400466 149614
rect 400702 149378 400874 149614
rect 400294 113934 400874 149378
rect 400294 113698 400466 113934
rect 400702 113698 400874 113934
rect 400294 113614 400874 113698
rect 400294 113378 400466 113614
rect 400702 113378 400874 113614
rect 400294 77934 400874 113378
rect 400294 77698 400466 77934
rect 400702 77698 400874 77934
rect 400294 77614 400874 77698
rect 400294 77378 400466 77614
rect 400702 77378 400874 77614
rect 400294 41934 400874 77378
rect 400294 41698 400466 41934
rect 400702 41698 400874 41934
rect 400294 41614 400874 41698
rect 400294 41378 400466 41614
rect 400702 41378 400874 41614
rect 400294 5934 400874 41378
rect 400294 5698 400466 5934
rect 400702 5698 400874 5934
rect 400294 5614 400874 5698
rect 400294 5378 400466 5614
rect 400702 5378 400874 5614
rect 400294 -2186 400874 5378
rect 400294 -2422 400466 -2186
rect 400702 -2422 400874 -2186
rect 400294 -2506 400874 -2422
rect 400294 -2742 400466 -2506
rect 400702 -2742 400874 -2506
rect 400294 -3674 400874 -2742
rect 403774 693414 404354 707962
rect 403774 693178 403946 693414
rect 404182 693178 404354 693414
rect 403774 693094 404354 693178
rect 403774 692858 403946 693094
rect 404182 692858 404354 693094
rect 403774 657414 404354 692858
rect 403774 657178 403946 657414
rect 404182 657178 404354 657414
rect 403774 657094 404354 657178
rect 403774 656858 403946 657094
rect 404182 656858 404354 657094
rect 403774 621414 404354 656858
rect 403774 621178 403946 621414
rect 404182 621178 404354 621414
rect 403774 621094 404354 621178
rect 403774 620858 403946 621094
rect 404182 620858 404354 621094
rect 403774 585414 404354 620858
rect 403774 585178 403946 585414
rect 404182 585178 404354 585414
rect 403774 585094 404354 585178
rect 403774 584858 403946 585094
rect 404182 584858 404354 585094
rect 403774 549414 404354 584858
rect 403774 549178 403946 549414
rect 404182 549178 404354 549414
rect 403774 549094 404354 549178
rect 403774 548858 403946 549094
rect 404182 548858 404354 549094
rect 403774 513414 404354 548858
rect 403774 513178 403946 513414
rect 404182 513178 404354 513414
rect 403774 513094 404354 513178
rect 403774 512858 403946 513094
rect 404182 512858 404354 513094
rect 403774 477414 404354 512858
rect 403774 477178 403946 477414
rect 404182 477178 404354 477414
rect 403774 477094 404354 477178
rect 403774 476858 403946 477094
rect 404182 476858 404354 477094
rect 403774 441414 404354 476858
rect 403774 441178 403946 441414
rect 404182 441178 404354 441414
rect 403774 441094 404354 441178
rect 403774 440858 403946 441094
rect 404182 440858 404354 441094
rect 403774 405414 404354 440858
rect 403774 405178 403946 405414
rect 404182 405178 404354 405414
rect 403774 405094 404354 405178
rect 403774 404858 403946 405094
rect 404182 404858 404354 405094
rect 403774 369414 404354 404858
rect 403774 369178 403946 369414
rect 404182 369178 404354 369414
rect 403774 369094 404354 369178
rect 403774 368858 403946 369094
rect 404182 368858 404354 369094
rect 403774 333414 404354 368858
rect 403774 333178 403946 333414
rect 404182 333178 404354 333414
rect 403774 333094 404354 333178
rect 403774 332858 403946 333094
rect 404182 332858 404354 333094
rect 403774 297414 404354 332858
rect 403774 297178 403946 297414
rect 404182 297178 404354 297414
rect 403774 297094 404354 297178
rect 403774 296858 403946 297094
rect 404182 296858 404354 297094
rect 403774 261414 404354 296858
rect 403774 261178 403946 261414
rect 404182 261178 404354 261414
rect 403774 261094 404354 261178
rect 403774 260858 403946 261094
rect 404182 260858 404354 261094
rect 403774 225414 404354 260858
rect 403774 225178 403946 225414
rect 404182 225178 404354 225414
rect 403774 225094 404354 225178
rect 403774 224858 403946 225094
rect 404182 224858 404354 225094
rect 403774 189414 404354 224858
rect 403774 189178 403946 189414
rect 404182 189178 404354 189414
rect 403774 189094 404354 189178
rect 403774 188858 403946 189094
rect 404182 188858 404354 189094
rect 403774 153414 404354 188858
rect 403774 153178 403946 153414
rect 404182 153178 404354 153414
rect 403774 153094 404354 153178
rect 403774 152858 403946 153094
rect 404182 152858 404354 153094
rect 403774 117414 404354 152858
rect 403774 117178 403946 117414
rect 404182 117178 404354 117414
rect 403774 117094 404354 117178
rect 403774 116858 403946 117094
rect 404182 116858 404354 117094
rect 403774 81414 404354 116858
rect 403774 81178 403946 81414
rect 404182 81178 404354 81414
rect 403774 81094 404354 81178
rect 403774 80858 403946 81094
rect 404182 80858 404354 81094
rect 403774 45414 404354 80858
rect 403774 45178 403946 45414
rect 404182 45178 404354 45414
rect 403774 45094 404354 45178
rect 403774 44858 403946 45094
rect 404182 44858 404354 45094
rect 403774 9414 404354 44858
rect 403774 9178 403946 9414
rect 404182 9178 404354 9414
rect 403774 9094 404354 9178
rect 403774 8858 403946 9094
rect 404182 8858 404354 9094
rect 403774 -4026 404354 8858
rect 403774 -4262 403946 -4026
rect 404182 -4262 404354 -4026
rect 403774 -4346 404354 -4262
rect 403774 -4582 403946 -4346
rect 404182 -4582 404354 -4346
rect 403774 -5514 404354 -4582
rect 407254 696894 407834 709802
rect 425254 711278 425834 711290
rect 425254 711042 425426 711278
rect 425662 711042 425834 711278
rect 425254 710958 425834 711042
rect 425254 710722 425426 710958
rect 425662 710722 425834 710958
rect 421774 709438 422354 709450
rect 421774 709202 421946 709438
rect 422182 709202 422354 709438
rect 421774 709118 422354 709202
rect 421774 708882 421946 709118
rect 422182 708882 422354 709118
rect 418294 707598 418874 707610
rect 418294 707362 418466 707598
rect 418702 707362 418874 707598
rect 418294 707278 418874 707362
rect 418294 707042 418466 707278
rect 418702 707042 418874 707278
rect 407254 696658 407426 696894
rect 407662 696658 407834 696894
rect 407254 696574 407834 696658
rect 407254 696338 407426 696574
rect 407662 696338 407834 696574
rect 407254 660894 407834 696338
rect 407254 660658 407426 660894
rect 407662 660658 407834 660894
rect 407254 660574 407834 660658
rect 407254 660338 407426 660574
rect 407662 660338 407834 660574
rect 407254 624894 407834 660338
rect 407254 624658 407426 624894
rect 407662 624658 407834 624894
rect 407254 624574 407834 624658
rect 407254 624338 407426 624574
rect 407662 624338 407834 624574
rect 407254 588894 407834 624338
rect 407254 588658 407426 588894
rect 407662 588658 407834 588894
rect 407254 588574 407834 588658
rect 407254 588338 407426 588574
rect 407662 588338 407834 588574
rect 407254 552894 407834 588338
rect 407254 552658 407426 552894
rect 407662 552658 407834 552894
rect 407254 552574 407834 552658
rect 407254 552338 407426 552574
rect 407662 552338 407834 552574
rect 407254 516894 407834 552338
rect 407254 516658 407426 516894
rect 407662 516658 407834 516894
rect 407254 516574 407834 516658
rect 407254 516338 407426 516574
rect 407662 516338 407834 516574
rect 407254 480894 407834 516338
rect 407254 480658 407426 480894
rect 407662 480658 407834 480894
rect 407254 480574 407834 480658
rect 407254 480338 407426 480574
rect 407662 480338 407834 480574
rect 407254 444894 407834 480338
rect 407254 444658 407426 444894
rect 407662 444658 407834 444894
rect 407254 444574 407834 444658
rect 407254 444338 407426 444574
rect 407662 444338 407834 444574
rect 407254 408894 407834 444338
rect 407254 408658 407426 408894
rect 407662 408658 407834 408894
rect 407254 408574 407834 408658
rect 407254 408338 407426 408574
rect 407662 408338 407834 408574
rect 407254 372894 407834 408338
rect 407254 372658 407426 372894
rect 407662 372658 407834 372894
rect 407254 372574 407834 372658
rect 407254 372338 407426 372574
rect 407662 372338 407834 372574
rect 407254 336894 407834 372338
rect 407254 336658 407426 336894
rect 407662 336658 407834 336894
rect 407254 336574 407834 336658
rect 407254 336338 407426 336574
rect 407662 336338 407834 336574
rect 407254 300894 407834 336338
rect 407254 300658 407426 300894
rect 407662 300658 407834 300894
rect 407254 300574 407834 300658
rect 407254 300338 407426 300574
rect 407662 300338 407834 300574
rect 407254 264894 407834 300338
rect 407254 264658 407426 264894
rect 407662 264658 407834 264894
rect 407254 264574 407834 264658
rect 407254 264338 407426 264574
rect 407662 264338 407834 264574
rect 407254 228894 407834 264338
rect 407254 228658 407426 228894
rect 407662 228658 407834 228894
rect 407254 228574 407834 228658
rect 407254 228338 407426 228574
rect 407662 228338 407834 228574
rect 407254 192894 407834 228338
rect 407254 192658 407426 192894
rect 407662 192658 407834 192894
rect 407254 192574 407834 192658
rect 407254 192338 407426 192574
rect 407662 192338 407834 192574
rect 407254 156894 407834 192338
rect 407254 156658 407426 156894
rect 407662 156658 407834 156894
rect 407254 156574 407834 156658
rect 407254 156338 407426 156574
rect 407662 156338 407834 156574
rect 407254 120894 407834 156338
rect 407254 120658 407426 120894
rect 407662 120658 407834 120894
rect 407254 120574 407834 120658
rect 407254 120338 407426 120574
rect 407662 120338 407834 120574
rect 407254 84894 407834 120338
rect 407254 84658 407426 84894
rect 407662 84658 407834 84894
rect 407254 84574 407834 84658
rect 407254 84338 407426 84574
rect 407662 84338 407834 84574
rect 407254 48894 407834 84338
rect 407254 48658 407426 48894
rect 407662 48658 407834 48894
rect 407254 48574 407834 48658
rect 407254 48338 407426 48574
rect 407662 48338 407834 48574
rect 407254 12894 407834 48338
rect 407254 12658 407426 12894
rect 407662 12658 407834 12894
rect 407254 12574 407834 12658
rect 407254 12338 407426 12574
rect 407662 12338 407834 12574
rect 389254 -7022 389426 -6786
rect 389662 -7022 389834 -6786
rect 389254 -7106 389834 -7022
rect 389254 -7342 389426 -7106
rect 389662 -7342 389834 -7106
rect 389254 -7354 389834 -7342
rect 407254 -5866 407834 12338
rect 414814 705758 415394 705770
rect 414814 705522 414986 705758
rect 415222 705522 415394 705758
rect 414814 705438 415394 705522
rect 414814 705202 414986 705438
rect 415222 705202 415394 705438
rect 414814 668454 415394 705202
rect 414814 668218 414986 668454
rect 415222 668218 415394 668454
rect 414814 668134 415394 668218
rect 414814 667898 414986 668134
rect 415222 667898 415394 668134
rect 414814 632454 415394 667898
rect 414814 632218 414986 632454
rect 415222 632218 415394 632454
rect 414814 632134 415394 632218
rect 414814 631898 414986 632134
rect 415222 631898 415394 632134
rect 414814 596454 415394 631898
rect 414814 596218 414986 596454
rect 415222 596218 415394 596454
rect 414814 596134 415394 596218
rect 414814 595898 414986 596134
rect 415222 595898 415394 596134
rect 414814 560454 415394 595898
rect 414814 560218 414986 560454
rect 415222 560218 415394 560454
rect 414814 560134 415394 560218
rect 414814 559898 414986 560134
rect 415222 559898 415394 560134
rect 414814 524454 415394 559898
rect 414814 524218 414986 524454
rect 415222 524218 415394 524454
rect 414814 524134 415394 524218
rect 414814 523898 414986 524134
rect 415222 523898 415394 524134
rect 414814 488454 415394 523898
rect 414814 488218 414986 488454
rect 415222 488218 415394 488454
rect 414814 488134 415394 488218
rect 414814 487898 414986 488134
rect 415222 487898 415394 488134
rect 414814 452454 415394 487898
rect 414814 452218 414986 452454
rect 415222 452218 415394 452454
rect 414814 452134 415394 452218
rect 414814 451898 414986 452134
rect 415222 451898 415394 452134
rect 414814 416454 415394 451898
rect 414814 416218 414986 416454
rect 415222 416218 415394 416454
rect 414814 416134 415394 416218
rect 414814 415898 414986 416134
rect 415222 415898 415394 416134
rect 414814 380454 415394 415898
rect 414814 380218 414986 380454
rect 415222 380218 415394 380454
rect 414814 380134 415394 380218
rect 414814 379898 414986 380134
rect 415222 379898 415394 380134
rect 414814 344454 415394 379898
rect 414814 344218 414986 344454
rect 415222 344218 415394 344454
rect 414814 344134 415394 344218
rect 414814 343898 414986 344134
rect 415222 343898 415394 344134
rect 414814 308454 415394 343898
rect 414814 308218 414986 308454
rect 415222 308218 415394 308454
rect 414814 308134 415394 308218
rect 414814 307898 414986 308134
rect 415222 307898 415394 308134
rect 414814 272454 415394 307898
rect 414814 272218 414986 272454
rect 415222 272218 415394 272454
rect 414814 272134 415394 272218
rect 414814 271898 414986 272134
rect 415222 271898 415394 272134
rect 414814 236454 415394 271898
rect 414814 236218 414986 236454
rect 415222 236218 415394 236454
rect 414814 236134 415394 236218
rect 414814 235898 414986 236134
rect 415222 235898 415394 236134
rect 414814 200454 415394 235898
rect 414814 200218 414986 200454
rect 415222 200218 415394 200454
rect 414814 200134 415394 200218
rect 414814 199898 414986 200134
rect 415222 199898 415394 200134
rect 414814 164454 415394 199898
rect 414814 164218 414986 164454
rect 415222 164218 415394 164454
rect 414814 164134 415394 164218
rect 414814 163898 414986 164134
rect 415222 163898 415394 164134
rect 414814 128454 415394 163898
rect 414814 128218 414986 128454
rect 415222 128218 415394 128454
rect 414814 128134 415394 128218
rect 414814 127898 414986 128134
rect 415222 127898 415394 128134
rect 414814 92454 415394 127898
rect 414814 92218 414986 92454
rect 415222 92218 415394 92454
rect 414814 92134 415394 92218
rect 414814 91898 414986 92134
rect 415222 91898 415394 92134
rect 414814 56454 415394 91898
rect 414814 56218 414986 56454
rect 415222 56218 415394 56454
rect 414814 56134 415394 56218
rect 414814 55898 414986 56134
rect 415222 55898 415394 56134
rect 414814 20454 415394 55898
rect 414814 20218 414986 20454
rect 415222 20218 415394 20454
rect 414814 20134 415394 20218
rect 414814 19898 414986 20134
rect 415222 19898 415394 20134
rect 414814 -1266 415394 19898
rect 414814 -1502 414986 -1266
rect 415222 -1502 415394 -1266
rect 414814 -1586 415394 -1502
rect 414814 -1822 414986 -1586
rect 415222 -1822 415394 -1586
rect 414814 -1834 415394 -1822
rect 418294 671934 418874 707042
rect 418294 671698 418466 671934
rect 418702 671698 418874 671934
rect 418294 671614 418874 671698
rect 418294 671378 418466 671614
rect 418702 671378 418874 671614
rect 418294 635934 418874 671378
rect 418294 635698 418466 635934
rect 418702 635698 418874 635934
rect 418294 635614 418874 635698
rect 418294 635378 418466 635614
rect 418702 635378 418874 635614
rect 418294 599934 418874 635378
rect 418294 599698 418466 599934
rect 418702 599698 418874 599934
rect 418294 599614 418874 599698
rect 418294 599378 418466 599614
rect 418702 599378 418874 599614
rect 418294 563934 418874 599378
rect 418294 563698 418466 563934
rect 418702 563698 418874 563934
rect 418294 563614 418874 563698
rect 418294 563378 418466 563614
rect 418702 563378 418874 563614
rect 418294 527934 418874 563378
rect 418294 527698 418466 527934
rect 418702 527698 418874 527934
rect 418294 527614 418874 527698
rect 418294 527378 418466 527614
rect 418702 527378 418874 527614
rect 418294 491934 418874 527378
rect 418294 491698 418466 491934
rect 418702 491698 418874 491934
rect 418294 491614 418874 491698
rect 418294 491378 418466 491614
rect 418702 491378 418874 491614
rect 418294 455934 418874 491378
rect 418294 455698 418466 455934
rect 418702 455698 418874 455934
rect 418294 455614 418874 455698
rect 418294 455378 418466 455614
rect 418702 455378 418874 455614
rect 418294 419934 418874 455378
rect 418294 419698 418466 419934
rect 418702 419698 418874 419934
rect 418294 419614 418874 419698
rect 418294 419378 418466 419614
rect 418702 419378 418874 419614
rect 418294 383934 418874 419378
rect 418294 383698 418466 383934
rect 418702 383698 418874 383934
rect 418294 383614 418874 383698
rect 418294 383378 418466 383614
rect 418702 383378 418874 383614
rect 418294 347934 418874 383378
rect 418294 347698 418466 347934
rect 418702 347698 418874 347934
rect 418294 347614 418874 347698
rect 418294 347378 418466 347614
rect 418702 347378 418874 347614
rect 418294 311934 418874 347378
rect 418294 311698 418466 311934
rect 418702 311698 418874 311934
rect 418294 311614 418874 311698
rect 418294 311378 418466 311614
rect 418702 311378 418874 311614
rect 418294 275934 418874 311378
rect 418294 275698 418466 275934
rect 418702 275698 418874 275934
rect 418294 275614 418874 275698
rect 418294 275378 418466 275614
rect 418702 275378 418874 275614
rect 418294 239934 418874 275378
rect 418294 239698 418466 239934
rect 418702 239698 418874 239934
rect 418294 239614 418874 239698
rect 418294 239378 418466 239614
rect 418702 239378 418874 239614
rect 418294 203934 418874 239378
rect 418294 203698 418466 203934
rect 418702 203698 418874 203934
rect 418294 203614 418874 203698
rect 418294 203378 418466 203614
rect 418702 203378 418874 203614
rect 418294 167934 418874 203378
rect 418294 167698 418466 167934
rect 418702 167698 418874 167934
rect 418294 167614 418874 167698
rect 418294 167378 418466 167614
rect 418702 167378 418874 167614
rect 418294 131934 418874 167378
rect 418294 131698 418466 131934
rect 418702 131698 418874 131934
rect 418294 131614 418874 131698
rect 418294 131378 418466 131614
rect 418702 131378 418874 131614
rect 418294 95934 418874 131378
rect 418294 95698 418466 95934
rect 418702 95698 418874 95934
rect 418294 95614 418874 95698
rect 418294 95378 418466 95614
rect 418702 95378 418874 95614
rect 418294 59934 418874 95378
rect 418294 59698 418466 59934
rect 418702 59698 418874 59934
rect 418294 59614 418874 59698
rect 418294 59378 418466 59614
rect 418702 59378 418874 59614
rect 418294 23934 418874 59378
rect 418294 23698 418466 23934
rect 418702 23698 418874 23934
rect 418294 23614 418874 23698
rect 418294 23378 418466 23614
rect 418702 23378 418874 23614
rect 418294 -3106 418874 23378
rect 418294 -3342 418466 -3106
rect 418702 -3342 418874 -3106
rect 418294 -3426 418874 -3342
rect 418294 -3662 418466 -3426
rect 418702 -3662 418874 -3426
rect 418294 -3674 418874 -3662
rect 421774 675414 422354 708882
rect 421774 675178 421946 675414
rect 422182 675178 422354 675414
rect 421774 675094 422354 675178
rect 421774 674858 421946 675094
rect 422182 674858 422354 675094
rect 421774 639414 422354 674858
rect 421774 639178 421946 639414
rect 422182 639178 422354 639414
rect 421774 639094 422354 639178
rect 421774 638858 421946 639094
rect 422182 638858 422354 639094
rect 421774 603414 422354 638858
rect 421774 603178 421946 603414
rect 422182 603178 422354 603414
rect 421774 603094 422354 603178
rect 421774 602858 421946 603094
rect 422182 602858 422354 603094
rect 421774 567414 422354 602858
rect 421774 567178 421946 567414
rect 422182 567178 422354 567414
rect 421774 567094 422354 567178
rect 421774 566858 421946 567094
rect 422182 566858 422354 567094
rect 421774 531414 422354 566858
rect 421774 531178 421946 531414
rect 422182 531178 422354 531414
rect 421774 531094 422354 531178
rect 421774 530858 421946 531094
rect 422182 530858 422354 531094
rect 421774 495414 422354 530858
rect 421774 495178 421946 495414
rect 422182 495178 422354 495414
rect 421774 495094 422354 495178
rect 421774 494858 421946 495094
rect 422182 494858 422354 495094
rect 421774 459414 422354 494858
rect 421774 459178 421946 459414
rect 422182 459178 422354 459414
rect 421774 459094 422354 459178
rect 421774 458858 421946 459094
rect 422182 458858 422354 459094
rect 421774 423414 422354 458858
rect 421774 423178 421946 423414
rect 422182 423178 422354 423414
rect 421774 423094 422354 423178
rect 421774 422858 421946 423094
rect 422182 422858 422354 423094
rect 421774 387414 422354 422858
rect 421774 387178 421946 387414
rect 422182 387178 422354 387414
rect 421774 387094 422354 387178
rect 421774 386858 421946 387094
rect 422182 386858 422354 387094
rect 421774 351414 422354 386858
rect 421774 351178 421946 351414
rect 422182 351178 422354 351414
rect 421774 351094 422354 351178
rect 421774 350858 421946 351094
rect 422182 350858 422354 351094
rect 421774 315414 422354 350858
rect 421774 315178 421946 315414
rect 422182 315178 422354 315414
rect 421774 315094 422354 315178
rect 421774 314858 421946 315094
rect 422182 314858 422354 315094
rect 421774 279414 422354 314858
rect 421774 279178 421946 279414
rect 422182 279178 422354 279414
rect 421774 279094 422354 279178
rect 421774 278858 421946 279094
rect 422182 278858 422354 279094
rect 421774 243414 422354 278858
rect 421774 243178 421946 243414
rect 422182 243178 422354 243414
rect 421774 243094 422354 243178
rect 421774 242858 421946 243094
rect 422182 242858 422354 243094
rect 421774 207414 422354 242858
rect 421774 207178 421946 207414
rect 422182 207178 422354 207414
rect 421774 207094 422354 207178
rect 421774 206858 421946 207094
rect 422182 206858 422354 207094
rect 421774 171414 422354 206858
rect 421774 171178 421946 171414
rect 422182 171178 422354 171414
rect 421774 171094 422354 171178
rect 421774 170858 421946 171094
rect 422182 170858 422354 171094
rect 421774 135414 422354 170858
rect 421774 135178 421946 135414
rect 422182 135178 422354 135414
rect 421774 135094 422354 135178
rect 421774 134858 421946 135094
rect 422182 134858 422354 135094
rect 421774 99414 422354 134858
rect 421774 99178 421946 99414
rect 422182 99178 422354 99414
rect 421774 99094 422354 99178
rect 421774 98858 421946 99094
rect 422182 98858 422354 99094
rect 421774 63414 422354 98858
rect 421774 63178 421946 63414
rect 422182 63178 422354 63414
rect 421774 63094 422354 63178
rect 421774 62858 421946 63094
rect 422182 62858 422354 63094
rect 421774 27414 422354 62858
rect 421774 27178 421946 27414
rect 422182 27178 422354 27414
rect 421774 27094 422354 27178
rect 421774 26858 421946 27094
rect 422182 26858 422354 27094
rect 421774 -4946 422354 26858
rect 421774 -5182 421946 -4946
rect 422182 -5182 422354 -4946
rect 421774 -5266 422354 -5182
rect 421774 -5502 421946 -5266
rect 422182 -5502 422354 -5266
rect 421774 -5514 422354 -5502
rect 425254 678894 425834 710722
rect 443254 710358 443834 711290
rect 443254 710122 443426 710358
rect 443662 710122 443834 710358
rect 443254 710038 443834 710122
rect 443254 709802 443426 710038
rect 443662 709802 443834 710038
rect 439774 708518 440354 709450
rect 439774 708282 439946 708518
rect 440182 708282 440354 708518
rect 439774 708198 440354 708282
rect 439774 707962 439946 708198
rect 440182 707962 440354 708198
rect 436294 706678 436874 707610
rect 436294 706442 436466 706678
rect 436702 706442 436874 706678
rect 436294 706358 436874 706442
rect 436294 706122 436466 706358
rect 436702 706122 436874 706358
rect 425254 678658 425426 678894
rect 425662 678658 425834 678894
rect 425254 678574 425834 678658
rect 425254 678338 425426 678574
rect 425662 678338 425834 678574
rect 425254 642894 425834 678338
rect 425254 642658 425426 642894
rect 425662 642658 425834 642894
rect 425254 642574 425834 642658
rect 425254 642338 425426 642574
rect 425662 642338 425834 642574
rect 425254 606894 425834 642338
rect 425254 606658 425426 606894
rect 425662 606658 425834 606894
rect 425254 606574 425834 606658
rect 425254 606338 425426 606574
rect 425662 606338 425834 606574
rect 425254 570894 425834 606338
rect 425254 570658 425426 570894
rect 425662 570658 425834 570894
rect 425254 570574 425834 570658
rect 425254 570338 425426 570574
rect 425662 570338 425834 570574
rect 425254 534894 425834 570338
rect 425254 534658 425426 534894
rect 425662 534658 425834 534894
rect 425254 534574 425834 534658
rect 425254 534338 425426 534574
rect 425662 534338 425834 534574
rect 425254 498894 425834 534338
rect 425254 498658 425426 498894
rect 425662 498658 425834 498894
rect 425254 498574 425834 498658
rect 425254 498338 425426 498574
rect 425662 498338 425834 498574
rect 425254 462894 425834 498338
rect 425254 462658 425426 462894
rect 425662 462658 425834 462894
rect 425254 462574 425834 462658
rect 425254 462338 425426 462574
rect 425662 462338 425834 462574
rect 425254 426894 425834 462338
rect 425254 426658 425426 426894
rect 425662 426658 425834 426894
rect 425254 426574 425834 426658
rect 425254 426338 425426 426574
rect 425662 426338 425834 426574
rect 425254 390894 425834 426338
rect 425254 390658 425426 390894
rect 425662 390658 425834 390894
rect 425254 390574 425834 390658
rect 425254 390338 425426 390574
rect 425662 390338 425834 390574
rect 425254 354894 425834 390338
rect 425254 354658 425426 354894
rect 425662 354658 425834 354894
rect 425254 354574 425834 354658
rect 425254 354338 425426 354574
rect 425662 354338 425834 354574
rect 425254 318894 425834 354338
rect 425254 318658 425426 318894
rect 425662 318658 425834 318894
rect 425254 318574 425834 318658
rect 425254 318338 425426 318574
rect 425662 318338 425834 318574
rect 425254 282894 425834 318338
rect 425254 282658 425426 282894
rect 425662 282658 425834 282894
rect 425254 282574 425834 282658
rect 425254 282338 425426 282574
rect 425662 282338 425834 282574
rect 425254 246894 425834 282338
rect 425254 246658 425426 246894
rect 425662 246658 425834 246894
rect 425254 246574 425834 246658
rect 425254 246338 425426 246574
rect 425662 246338 425834 246574
rect 425254 210894 425834 246338
rect 425254 210658 425426 210894
rect 425662 210658 425834 210894
rect 425254 210574 425834 210658
rect 425254 210338 425426 210574
rect 425662 210338 425834 210574
rect 425254 174894 425834 210338
rect 425254 174658 425426 174894
rect 425662 174658 425834 174894
rect 425254 174574 425834 174658
rect 425254 174338 425426 174574
rect 425662 174338 425834 174574
rect 425254 138894 425834 174338
rect 425254 138658 425426 138894
rect 425662 138658 425834 138894
rect 425254 138574 425834 138658
rect 425254 138338 425426 138574
rect 425662 138338 425834 138574
rect 425254 102894 425834 138338
rect 425254 102658 425426 102894
rect 425662 102658 425834 102894
rect 425254 102574 425834 102658
rect 425254 102338 425426 102574
rect 425662 102338 425834 102574
rect 425254 66894 425834 102338
rect 425254 66658 425426 66894
rect 425662 66658 425834 66894
rect 425254 66574 425834 66658
rect 425254 66338 425426 66574
rect 425662 66338 425834 66574
rect 425254 30894 425834 66338
rect 425254 30658 425426 30894
rect 425662 30658 425834 30894
rect 425254 30574 425834 30658
rect 425254 30338 425426 30574
rect 425662 30338 425834 30574
rect 407254 -6102 407426 -5866
rect 407662 -6102 407834 -5866
rect 407254 -6186 407834 -6102
rect 407254 -6422 407426 -6186
rect 407662 -6422 407834 -6186
rect 407254 -7354 407834 -6422
rect 425254 -6786 425834 30338
rect 432814 704838 433394 705770
rect 432814 704602 432986 704838
rect 433222 704602 433394 704838
rect 432814 704518 433394 704602
rect 432814 704282 432986 704518
rect 433222 704282 433394 704518
rect 432814 686454 433394 704282
rect 432814 686218 432986 686454
rect 433222 686218 433394 686454
rect 432814 686134 433394 686218
rect 432814 685898 432986 686134
rect 433222 685898 433394 686134
rect 432814 650454 433394 685898
rect 432814 650218 432986 650454
rect 433222 650218 433394 650454
rect 432814 650134 433394 650218
rect 432814 649898 432986 650134
rect 433222 649898 433394 650134
rect 432814 614454 433394 649898
rect 432814 614218 432986 614454
rect 433222 614218 433394 614454
rect 432814 614134 433394 614218
rect 432814 613898 432986 614134
rect 433222 613898 433394 614134
rect 432814 578454 433394 613898
rect 432814 578218 432986 578454
rect 433222 578218 433394 578454
rect 432814 578134 433394 578218
rect 432814 577898 432986 578134
rect 433222 577898 433394 578134
rect 432814 542454 433394 577898
rect 432814 542218 432986 542454
rect 433222 542218 433394 542454
rect 432814 542134 433394 542218
rect 432814 541898 432986 542134
rect 433222 541898 433394 542134
rect 432814 506454 433394 541898
rect 432814 506218 432986 506454
rect 433222 506218 433394 506454
rect 432814 506134 433394 506218
rect 432814 505898 432986 506134
rect 433222 505898 433394 506134
rect 432814 470454 433394 505898
rect 432814 470218 432986 470454
rect 433222 470218 433394 470454
rect 432814 470134 433394 470218
rect 432814 469898 432986 470134
rect 433222 469898 433394 470134
rect 432814 434454 433394 469898
rect 432814 434218 432986 434454
rect 433222 434218 433394 434454
rect 432814 434134 433394 434218
rect 432814 433898 432986 434134
rect 433222 433898 433394 434134
rect 432814 398454 433394 433898
rect 432814 398218 432986 398454
rect 433222 398218 433394 398454
rect 432814 398134 433394 398218
rect 432814 397898 432986 398134
rect 433222 397898 433394 398134
rect 432814 362454 433394 397898
rect 432814 362218 432986 362454
rect 433222 362218 433394 362454
rect 432814 362134 433394 362218
rect 432814 361898 432986 362134
rect 433222 361898 433394 362134
rect 432814 326454 433394 361898
rect 432814 326218 432986 326454
rect 433222 326218 433394 326454
rect 432814 326134 433394 326218
rect 432814 325898 432986 326134
rect 433222 325898 433394 326134
rect 432814 290454 433394 325898
rect 432814 290218 432986 290454
rect 433222 290218 433394 290454
rect 432814 290134 433394 290218
rect 432814 289898 432986 290134
rect 433222 289898 433394 290134
rect 432814 254454 433394 289898
rect 432814 254218 432986 254454
rect 433222 254218 433394 254454
rect 432814 254134 433394 254218
rect 432814 253898 432986 254134
rect 433222 253898 433394 254134
rect 432814 218454 433394 253898
rect 432814 218218 432986 218454
rect 433222 218218 433394 218454
rect 432814 218134 433394 218218
rect 432814 217898 432986 218134
rect 433222 217898 433394 218134
rect 432814 182454 433394 217898
rect 432814 182218 432986 182454
rect 433222 182218 433394 182454
rect 432814 182134 433394 182218
rect 432814 181898 432986 182134
rect 433222 181898 433394 182134
rect 432814 146454 433394 181898
rect 432814 146218 432986 146454
rect 433222 146218 433394 146454
rect 432814 146134 433394 146218
rect 432814 145898 432986 146134
rect 433222 145898 433394 146134
rect 432814 110454 433394 145898
rect 432814 110218 432986 110454
rect 433222 110218 433394 110454
rect 432814 110134 433394 110218
rect 432814 109898 432986 110134
rect 433222 109898 433394 110134
rect 432814 74454 433394 109898
rect 432814 74218 432986 74454
rect 433222 74218 433394 74454
rect 432814 74134 433394 74218
rect 432814 73898 432986 74134
rect 433222 73898 433394 74134
rect 432814 38454 433394 73898
rect 432814 38218 432986 38454
rect 433222 38218 433394 38454
rect 432814 38134 433394 38218
rect 432814 37898 432986 38134
rect 433222 37898 433394 38134
rect 432814 2454 433394 37898
rect 432814 2218 432986 2454
rect 433222 2218 433394 2454
rect 432814 2134 433394 2218
rect 432814 1898 432986 2134
rect 433222 1898 433394 2134
rect 432814 -346 433394 1898
rect 432814 -582 432986 -346
rect 433222 -582 433394 -346
rect 432814 -666 433394 -582
rect 432814 -902 432986 -666
rect 433222 -902 433394 -666
rect 432814 -1834 433394 -902
rect 436294 689934 436874 706122
rect 436294 689698 436466 689934
rect 436702 689698 436874 689934
rect 436294 689614 436874 689698
rect 436294 689378 436466 689614
rect 436702 689378 436874 689614
rect 436294 653934 436874 689378
rect 436294 653698 436466 653934
rect 436702 653698 436874 653934
rect 436294 653614 436874 653698
rect 436294 653378 436466 653614
rect 436702 653378 436874 653614
rect 436294 617934 436874 653378
rect 436294 617698 436466 617934
rect 436702 617698 436874 617934
rect 436294 617614 436874 617698
rect 436294 617378 436466 617614
rect 436702 617378 436874 617614
rect 436294 581934 436874 617378
rect 436294 581698 436466 581934
rect 436702 581698 436874 581934
rect 436294 581614 436874 581698
rect 436294 581378 436466 581614
rect 436702 581378 436874 581614
rect 436294 545934 436874 581378
rect 436294 545698 436466 545934
rect 436702 545698 436874 545934
rect 436294 545614 436874 545698
rect 436294 545378 436466 545614
rect 436702 545378 436874 545614
rect 436294 509934 436874 545378
rect 436294 509698 436466 509934
rect 436702 509698 436874 509934
rect 436294 509614 436874 509698
rect 436294 509378 436466 509614
rect 436702 509378 436874 509614
rect 436294 473934 436874 509378
rect 436294 473698 436466 473934
rect 436702 473698 436874 473934
rect 436294 473614 436874 473698
rect 436294 473378 436466 473614
rect 436702 473378 436874 473614
rect 436294 437934 436874 473378
rect 436294 437698 436466 437934
rect 436702 437698 436874 437934
rect 436294 437614 436874 437698
rect 436294 437378 436466 437614
rect 436702 437378 436874 437614
rect 436294 401934 436874 437378
rect 436294 401698 436466 401934
rect 436702 401698 436874 401934
rect 436294 401614 436874 401698
rect 436294 401378 436466 401614
rect 436702 401378 436874 401614
rect 436294 365934 436874 401378
rect 436294 365698 436466 365934
rect 436702 365698 436874 365934
rect 436294 365614 436874 365698
rect 436294 365378 436466 365614
rect 436702 365378 436874 365614
rect 436294 329934 436874 365378
rect 436294 329698 436466 329934
rect 436702 329698 436874 329934
rect 436294 329614 436874 329698
rect 436294 329378 436466 329614
rect 436702 329378 436874 329614
rect 436294 293934 436874 329378
rect 436294 293698 436466 293934
rect 436702 293698 436874 293934
rect 436294 293614 436874 293698
rect 436294 293378 436466 293614
rect 436702 293378 436874 293614
rect 436294 257934 436874 293378
rect 436294 257698 436466 257934
rect 436702 257698 436874 257934
rect 436294 257614 436874 257698
rect 436294 257378 436466 257614
rect 436702 257378 436874 257614
rect 436294 221934 436874 257378
rect 436294 221698 436466 221934
rect 436702 221698 436874 221934
rect 436294 221614 436874 221698
rect 436294 221378 436466 221614
rect 436702 221378 436874 221614
rect 436294 185934 436874 221378
rect 436294 185698 436466 185934
rect 436702 185698 436874 185934
rect 436294 185614 436874 185698
rect 436294 185378 436466 185614
rect 436702 185378 436874 185614
rect 436294 149934 436874 185378
rect 436294 149698 436466 149934
rect 436702 149698 436874 149934
rect 436294 149614 436874 149698
rect 436294 149378 436466 149614
rect 436702 149378 436874 149614
rect 436294 113934 436874 149378
rect 436294 113698 436466 113934
rect 436702 113698 436874 113934
rect 436294 113614 436874 113698
rect 436294 113378 436466 113614
rect 436702 113378 436874 113614
rect 436294 77934 436874 113378
rect 436294 77698 436466 77934
rect 436702 77698 436874 77934
rect 436294 77614 436874 77698
rect 436294 77378 436466 77614
rect 436702 77378 436874 77614
rect 436294 41934 436874 77378
rect 436294 41698 436466 41934
rect 436702 41698 436874 41934
rect 436294 41614 436874 41698
rect 436294 41378 436466 41614
rect 436702 41378 436874 41614
rect 436294 5934 436874 41378
rect 436294 5698 436466 5934
rect 436702 5698 436874 5934
rect 436294 5614 436874 5698
rect 436294 5378 436466 5614
rect 436702 5378 436874 5614
rect 436294 -2186 436874 5378
rect 436294 -2422 436466 -2186
rect 436702 -2422 436874 -2186
rect 436294 -2506 436874 -2422
rect 436294 -2742 436466 -2506
rect 436702 -2742 436874 -2506
rect 436294 -3674 436874 -2742
rect 439774 693414 440354 707962
rect 439774 693178 439946 693414
rect 440182 693178 440354 693414
rect 439774 693094 440354 693178
rect 439774 692858 439946 693094
rect 440182 692858 440354 693094
rect 439774 657414 440354 692858
rect 439774 657178 439946 657414
rect 440182 657178 440354 657414
rect 439774 657094 440354 657178
rect 439774 656858 439946 657094
rect 440182 656858 440354 657094
rect 439774 621414 440354 656858
rect 439774 621178 439946 621414
rect 440182 621178 440354 621414
rect 439774 621094 440354 621178
rect 439774 620858 439946 621094
rect 440182 620858 440354 621094
rect 439774 585414 440354 620858
rect 439774 585178 439946 585414
rect 440182 585178 440354 585414
rect 439774 585094 440354 585178
rect 439774 584858 439946 585094
rect 440182 584858 440354 585094
rect 439774 549414 440354 584858
rect 439774 549178 439946 549414
rect 440182 549178 440354 549414
rect 439774 549094 440354 549178
rect 439774 548858 439946 549094
rect 440182 548858 440354 549094
rect 439774 513414 440354 548858
rect 439774 513178 439946 513414
rect 440182 513178 440354 513414
rect 439774 513094 440354 513178
rect 439774 512858 439946 513094
rect 440182 512858 440354 513094
rect 439774 477414 440354 512858
rect 439774 477178 439946 477414
rect 440182 477178 440354 477414
rect 439774 477094 440354 477178
rect 439774 476858 439946 477094
rect 440182 476858 440354 477094
rect 439774 441414 440354 476858
rect 439774 441178 439946 441414
rect 440182 441178 440354 441414
rect 439774 441094 440354 441178
rect 439774 440858 439946 441094
rect 440182 440858 440354 441094
rect 439774 405414 440354 440858
rect 439774 405178 439946 405414
rect 440182 405178 440354 405414
rect 439774 405094 440354 405178
rect 439774 404858 439946 405094
rect 440182 404858 440354 405094
rect 439774 369414 440354 404858
rect 439774 369178 439946 369414
rect 440182 369178 440354 369414
rect 439774 369094 440354 369178
rect 439774 368858 439946 369094
rect 440182 368858 440354 369094
rect 439774 333414 440354 368858
rect 439774 333178 439946 333414
rect 440182 333178 440354 333414
rect 439774 333094 440354 333178
rect 439774 332858 439946 333094
rect 440182 332858 440354 333094
rect 439774 297414 440354 332858
rect 439774 297178 439946 297414
rect 440182 297178 440354 297414
rect 439774 297094 440354 297178
rect 439774 296858 439946 297094
rect 440182 296858 440354 297094
rect 439774 261414 440354 296858
rect 439774 261178 439946 261414
rect 440182 261178 440354 261414
rect 439774 261094 440354 261178
rect 439774 260858 439946 261094
rect 440182 260858 440354 261094
rect 439774 225414 440354 260858
rect 439774 225178 439946 225414
rect 440182 225178 440354 225414
rect 439774 225094 440354 225178
rect 439774 224858 439946 225094
rect 440182 224858 440354 225094
rect 439774 189414 440354 224858
rect 439774 189178 439946 189414
rect 440182 189178 440354 189414
rect 439774 189094 440354 189178
rect 439774 188858 439946 189094
rect 440182 188858 440354 189094
rect 439774 153414 440354 188858
rect 439774 153178 439946 153414
rect 440182 153178 440354 153414
rect 439774 153094 440354 153178
rect 439774 152858 439946 153094
rect 440182 152858 440354 153094
rect 439774 117414 440354 152858
rect 439774 117178 439946 117414
rect 440182 117178 440354 117414
rect 439774 117094 440354 117178
rect 439774 116858 439946 117094
rect 440182 116858 440354 117094
rect 439774 81414 440354 116858
rect 439774 81178 439946 81414
rect 440182 81178 440354 81414
rect 439774 81094 440354 81178
rect 439774 80858 439946 81094
rect 440182 80858 440354 81094
rect 439774 45414 440354 80858
rect 439774 45178 439946 45414
rect 440182 45178 440354 45414
rect 439774 45094 440354 45178
rect 439774 44858 439946 45094
rect 440182 44858 440354 45094
rect 439774 9414 440354 44858
rect 439774 9178 439946 9414
rect 440182 9178 440354 9414
rect 439774 9094 440354 9178
rect 439774 8858 439946 9094
rect 440182 8858 440354 9094
rect 439774 -4026 440354 8858
rect 439774 -4262 439946 -4026
rect 440182 -4262 440354 -4026
rect 439774 -4346 440354 -4262
rect 439774 -4582 439946 -4346
rect 440182 -4582 440354 -4346
rect 439774 -5514 440354 -4582
rect 443254 696894 443834 709802
rect 461254 711278 461834 711290
rect 461254 711042 461426 711278
rect 461662 711042 461834 711278
rect 461254 710958 461834 711042
rect 461254 710722 461426 710958
rect 461662 710722 461834 710958
rect 457774 709438 458354 709450
rect 457774 709202 457946 709438
rect 458182 709202 458354 709438
rect 457774 709118 458354 709202
rect 457774 708882 457946 709118
rect 458182 708882 458354 709118
rect 454294 707598 454874 707610
rect 454294 707362 454466 707598
rect 454702 707362 454874 707598
rect 454294 707278 454874 707362
rect 454294 707042 454466 707278
rect 454702 707042 454874 707278
rect 443254 696658 443426 696894
rect 443662 696658 443834 696894
rect 443254 696574 443834 696658
rect 443254 696338 443426 696574
rect 443662 696338 443834 696574
rect 443254 660894 443834 696338
rect 443254 660658 443426 660894
rect 443662 660658 443834 660894
rect 443254 660574 443834 660658
rect 443254 660338 443426 660574
rect 443662 660338 443834 660574
rect 443254 624894 443834 660338
rect 443254 624658 443426 624894
rect 443662 624658 443834 624894
rect 443254 624574 443834 624658
rect 443254 624338 443426 624574
rect 443662 624338 443834 624574
rect 443254 588894 443834 624338
rect 443254 588658 443426 588894
rect 443662 588658 443834 588894
rect 443254 588574 443834 588658
rect 443254 588338 443426 588574
rect 443662 588338 443834 588574
rect 443254 552894 443834 588338
rect 443254 552658 443426 552894
rect 443662 552658 443834 552894
rect 443254 552574 443834 552658
rect 443254 552338 443426 552574
rect 443662 552338 443834 552574
rect 443254 516894 443834 552338
rect 443254 516658 443426 516894
rect 443662 516658 443834 516894
rect 443254 516574 443834 516658
rect 443254 516338 443426 516574
rect 443662 516338 443834 516574
rect 443254 480894 443834 516338
rect 443254 480658 443426 480894
rect 443662 480658 443834 480894
rect 443254 480574 443834 480658
rect 443254 480338 443426 480574
rect 443662 480338 443834 480574
rect 443254 444894 443834 480338
rect 443254 444658 443426 444894
rect 443662 444658 443834 444894
rect 443254 444574 443834 444658
rect 443254 444338 443426 444574
rect 443662 444338 443834 444574
rect 443254 408894 443834 444338
rect 443254 408658 443426 408894
rect 443662 408658 443834 408894
rect 443254 408574 443834 408658
rect 443254 408338 443426 408574
rect 443662 408338 443834 408574
rect 443254 372894 443834 408338
rect 443254 372658 443426 372894
rect 443662 372658 443834 372894
rect 443254 372574 443834 372658
rect 443254 372338 443426 372574
rect 443662 372338 443834 372574
rect 443254 336894 443834 372338
rect 443254 336658 443426 336894
rect 443662 336658 443834 336894
rect 443254 336574 443834 336658
rect 443254 336338 443426 336574
rect 443662 336338 443834 336574
rect 443254 300894 443834 336338
rect 443254 300658 443426 300894
rect 443662 300658 443834 300894
rect 443254 300574 443834 300658
rect 443254 300338 443426 300574
rect 443662 300338 443834 300574
rect 443254 264894 443834 300338
rect 443254 264658 443426 264894
rect 443662 264658 443834 264894
rect 443254 264574 443834 264658
rect 443254 264338 443426 264574
rect 443662 264338 443834 264574
rect 443254 228894 443834 264338
rect 443254 228658 443426 228894
rect 443662 228658 443834 228894
rect 443254 228574 443834 228658
rect 443254 228338 443426 228574
rect 443662 228338 443834 228574
rect 443254 192894 443834 228338
rect 443254 192658 443426 192894
rect 443662 192658 443834 192894
rect 443254 192574 443834 192658
rect 443254 192338 443426 192574
rect 443662 192338 443834 192574
rect 443254 156894 443834 192338
rect 443254 156658 443426 156894
rect 443662 156658 443834 156894
rect 443254 156574 443834 156658
rect 443254 156338 443426 156574
rect 443662 156338 443834 156574
rect 443254 120894 443834 156338
rect 443254 120658 443426 120894
rect 443662 120658 443834 120894
rect 443254 120574 443834 120658
rect 443254 120338 443426 120574
rect 443662 120338 443834 120574
rect 443254 84894 443834 120338
rect 443254 84658 443426 84894
rect 443662 84658 443834 84894
rect 443254 84574 443834 84658
rect 443254 84338 443426 84574
rect 443662 84338 443834 84574
rect 443254 48894 443834 84338
rect 443254 48658 443426 48894
rect 443662 48658 443834 48894
rect 443254 48574 443834 48658
rect 443254 48338 443426 48574
rect 443662 48338 443834 48574
rect 443254 12894 443834 48338
rect 443254 12658 443426 12894
rect 443662 12658 443834 12894
rect 443254 12574 443834 12658
rect 443254 12338 443426 12574
rect 443662 12338 443834 12574
rect 425254 -7022 425426 -6786
rect 425662 -7022 425834 -6786
rect 425254 -7106 425834 -7022
rect 425254 -7342 425426 -7106
rect 425662 -7342 425834 -7106
rect 425254 -7354 425834 -7342
rect 443254 -5866 443834 12338
rect 450814 705758 451394 705770
rect 450814 705522 450986 705758
rect 451222 705522 451394 705758
rect 450814 705438 451394 705522
rect 450814 705202 450986 705438
rect 451222 705202 451394 705438
rect 450814 668454 451394 705202
rect 450814 668218 450986 668454
rect 451222 668218 451394 668454
rect 450814 668134 451394 668218
rect 450814 667898 450986 668134
rect 451222 667898 451394 668134
rect 450814 632454 451394 667898
rect 450814 632218 450986 632454
rect 451222 632218 451394 632454
rect 450814 632134 451394 632218
rect 450814 631898 450986 632134
rect 451222 631898 451394 632134
rect 450814 596454 451394 631898
rect 450814 596218 450986 596454
rect 451222 596218 451394 596454
rect 450814 596134 451394 596218
rect 450814 595898 450986 596134
rect 451222 595898 451394 596134
rect 450814 560454 451394 595898
rect 450814 560218 450986 560454
rect 451222 560218 451394 560454
rect 450814 560134 451394 560218
rect 450814 559898 450986 560134
rect 451222 559898 451394 560134
rect 450814 524454 451394 559898
rect 450814 524218 450986 524454
rect 451222 524218 451394 524454
rect 450814 524134 451394 524218
rect 450814 523898 450986 524134
rect 451222 523898 451394 524134
rect 450814 488454 451394 523898
rect 450814 488218 450986 488454
rect 451222 488218 451394 488454
rect 450814 488134 451394 488218
rect 450814 487898 450986 488134
rect 451222 487898 451394 488134
rect 450814 452454 451394 487898
rect 450814 452218 450986 452454
rect 451222 452218 451394 452454
rect 450814 452134 451394 452218
rect 450814 451898 450986 452134
rect 451222 451898 451394 452134
rect 450814 416454 451394 451898
rect 450814 416218 450986 416454
rect 451222 416218 451394 416454
rect 450814 416134 451394 416218
rect 450814 415898 450986 416134
rect 451222 415898 451394 416134
rect 450814 380454 451394 415898
rect 450814 380218 450986 380454
rect 451222 380218 451394 380454
rect 450814 380134 451394 380218
rect 450814 379898 450986 380134
rect 451222 379898 451394 380134
rect 450814 344454 451394 379898
rect 450814 344218 450986 344454
rect 451222 344218 451394 344454
rect 450814 344134 451394 344218
rect 450814 343898 450986 344134
rect 451222 343898 451394 344134
rect 450814 308454 451394 343898
rect 450814 308218 450986 308454
rect 451222 308218 451394 308454
rect 450814 308134 451394 308218
rect 450814 307898 450986 308134
rect 451222 307898 451394 308134
rect 450814 272454 451394 307898
rect 450814 272218 450986 272454
rect 451222 272218 451394 272454
rect 450814 272134 451394 272218
rect 450814 271898 450986 272134
rect 451222 271898 451394 272134
rect 450814 236454 451394 271898
rect 450814 236218 450986 236454
rect 451222 236218 451394 236454
rect 450814 236134 451394 236218
rect 450814 235898 450986 236134
rect 451222 235898 451394 236134
rect 450814 200454 451394 235898
rect 450814 200218 450986 200454
rect 451222 200218 451394 200454
rect 450814 200134 451394 200218
rect 450814 199898 450986 200134
rect 451222 199898 451394 200134
rect 450814 164454 451394 199898
rect 450814 164218 450986 164454
rect 451222 164218 451394 164454
rect 450814 164134 451394 164218
rect 450814 163898 450986 164134
rect 451222 163898 451394 164134
rect 450814 128454 451394 163898
rect 450814 128218 450986 128454
rect 451222 128218 451394 128454
rect 450814 128134 451394 128218
rect 450814 127898 450986 128134
rect 451222 127898 451394 128134
rect 450814 92454 451394 127898
rect 450814 92218 450986 92454
rect 451222 92218 451394 92454
rect 450814 92134 451394 92218
rect 450814 91898 450986 92134
rect 451222 91898 451394 92134
rect 450814 56454 451394 91898
rect 450814 56218 450986 56454
rect 451222 56218 451394 56454
rect 450814 56134 451394 56218
rect 450814 55898 450986 56134
rect 451222 55898 451394 56134
rect 450814 20454 451394 55898
rect 450814 20218 450986 20454
rect 451222 20218 451394 20454
rect 450814 20134 451394 20218
rect 450814 19898 450986 20134
rect 451222 19898 451394 20134
rect 450814 -1266 451394 19898
rect 450814 -1502 450986 -1266
rect 451222 -1502 451394 -1266
rect 450814 -1586 451394 -1502
rect 450814 -1822 450986 -1586
rect 451222 -1822 451394 -1586
rect 450814 -1834 451394 -1822
rect 454294 671934 454874 707042
rect 454294 671698 454466 671934
rect 454702 671698 454874 671934
rect 454294 671614 454874 671698
rect 454294 671378 454466 671614
rect 454702 671378 454874 671614
rect 454294 635934 454874 671378
rect 454294 635698 454466 635934
rect 454702 635698 454874 635934
rect 454294 635614 454874 635698
rect 454294 635378 454466 635614
rect 454702 635378 454874 635614
rect 454294 599934 454874 635378
rect 454294 599698 454466 599934
rect 454702 599698 454874 599934
rect 454294 599614 454874 599698
rect 454294 599378 454466 599614
rect 454702 599378 454874 599614
rect 454294 563934 454874 599378
rect 454294 563698 454466 563934
rect 454702 563698 454874 563934
rect 454294 563614 454874 563698
rect 454294 563378 454466 563614
rect 454702 563378 454874 563614
rect 454294 527934 454874 563378
rect 454294 527698 454466 527934
rect 454702 527698 454874 527934
rect 454294 527614 454874 527698
rect 454294 527378 454466 527614
rect 454702 527378 454874 527614
rect 454294 491934 454874 527378
rect 454294 491698 454466 491934
rect 454702 491698 454874 491934
rect 454294 491614 454874 491698
rect 454294 491378 454466 491614
rect 454702 491378 454874 491614
rect 454294 455934 454874 491378
rect 454294 455698 454466 455934
rect 454702 455698 454874 455934
rect 454294 455614 454874 455698
rect 454294 455378 454466 455614
rect 454702 455378 454874 455614
rect 454294 419934 454874 455378
rect 454294 419698 454466 419934
rect 454702 419698 454874 419934
rect 454294 419614 454874 419698
rect 454294 419378 454466 419614
rect 454702 419378 454874 419614
rect 454294 383934 454874 419378
rect 454294 383698 454466 383934
rect 454702 383698 454874 383934
rect 454294 383614 454874 383698
rect 454294 383378 454466 383614
rect 454702 383378 454874 383614
rect 454294 347934 454874 383378
rect 454294 347698 454466 347934
rect 454702 347698 454874 347934
rect 454294 347614 454874 347698
rect 454294 347378 454466 347614
rect 454702 347378 454874 347614
rect 454294 311934 454874 347378
rect 454294 311698 454466 311934
rect 454702 311698 454874 311934
rect 454294 311614 454874 311698
rect 454294 311378 454466 311614
rect 454702 311378 454874 311614
rect 454294 275934 454874 311378
rect 454294 275698 454466 275934
rect 454702 275698 454874 275934
rect 454294 275614 454874 275698
rect 454294 275378 454466 275614
rect 454702 275378 454874 275614
rect 454294 239934 454874 275378
rect 454294 239698 454466 239934
rect 454702 239698 454874 239934
rect 454294 239614 454874 239698
rect 454294 239378 454466 239614
rect 454702 239378 454874 239614
rect 454294 203934 454874 239378
rect 454294 203698 454466 203934
rect 454702 203698 454874 203934
rect 454294 203614 454874 203698
rect 454294 203378 454466 203614
rect 454702 203378 454874 203614
rect 454294 167934 454874 203378
rect 454294 167698 454466 167934
rect 454702 167698 454874 167934
rect 454294 167614 454874 167698
rect 454294 167378 454466 167614
rect 454702 167378 454874 167614
rect 454294 131934 454874 167378
rect 454294 131698 454466 131934
rect 454702 131698 454874 131934
rect 454294 131614 454874 131698
rect 454294 131378 454466 131614
rect 454702 131378 454874 131614
rect 454294 95934 454874 131378
rect 454294 95698 454466 95934
rect 454702 95698 454874 95934
rect 454294 95614 454874 95698
rect 454294 95378 454466 95614
rect 454702 95378 454874 95614
rect 454294 59934 454874 95378
rect 454294 59698 454466 59934
rect 454702 59698 454874 59934
rect 454294 59614 454874 59698
rect 454294 59378 454466 59614
rect 454702 59378 454874 59614
rect 454294 23934 454874 59378
rect 454294 23698 454466 23934
rect 454702 23698 454874 23934
rect 454294 23614 454874 23698
rect 454294 23378 454466 23614
rect 454702 23378 454874 23614
rect 454294 -3106 454874 23378
rect 454294 -3342 454466 -3106
rect 454702 -3342 454874 -3106
rect 454294 -3426 454874 -3342
rect 454294 -3662 454466 -3426
rect 454702 -3662 454874 -3426
rect 454294 -3674 454874 -3662
rect 457774 675414 458354 708882
rect 457774 675178 457946 675414
rect 458182 675178 458354 675414
rect 457774 675094 458354 675178
rect 457774 674858 457946 675094
rect 458182 674858 458354 675094
rect 457774 639414 458354 674858
rect 457774 639178 457946 639414
rect 458182 639178 458354 639414
rect 457774 639094 458354 639178
rect 457774 638858 457946 639094
rect 458182 638858 458354 639094
rect 457774 603414 458354 638858
rect 457774 603178 457946 603414
rect 458182 603178 458354 603414
rect 457774 603094 458354 603178
rect 457774 602858 457946 603094
rect 458182 602858 458354 603094
rect 457774 567414 458354 602858
rect 457774 567178 457946 567414
rect 458182 567178 458354 567414
rect 457774 567094 458354 567178
rect 457774 566858 457946 567094
rect 458182 566858 458354 567094
rect 457774 531414 458354 566858
rect 457774 531178 457946 531414
rect 458182 531178 458354 531414
rect 457774 531094 458354 531178
rect 457774 530858 457946 531094
rect 458182 530858 458354 531094
rect 457774 495414 458354 530858
rect 457774 495178 457946 495414
rect 458182 495178 458354 495414
rect 457774 495094 458354 495178
rect 457774 494858 457946 495094
rect 458182 494858 458354 495094
rect 457774 459414 458354 494858
rect 457774 459178 457946 459414
rect 458182 459178 458354 459414
rect 457774 459094 458354 459178
rect 457774 458858 457946 459094
rect 458182 458858 458354 459094
rect 457774 423414 458354 458858
rect 457774 423178 457946 423414
rect 458182 423178 458354 423414
rect 457774 423094 458354 423178
rect 457774 422858 457946 423094
rect 458182 422858 458354 423094
rect 457774 387414 458354 422858
rect 457774 387178 457946 387414
rect 458182 387178 458354 387414
rect 457774 387094 458354 387178
rect 457774 386858 457946 387094
rect 458182 386858 458354 387094
rect 457774 351414 458354 386858
rect 457774 351178 457946 351414
rect 458182 351178 458354 351414
rect 457774 351094 458354 351178
rect 457774 350858 457946 351094
rect 458182 350858 458354 351094
rect 457774 315414 458354 350858
rect 457774 315178 457946 315414
rect 458182 315178 458354 315414
rect 457774 315094 458354 315178
rect 457774 314858 457946 315094
rect 458182 314858 458354 315094
rect 457774 279414 458354 314858
rect 457774 279178 457946 279414
rect 458182 279178 458354 279414
rect 457774 279094 458354 279178
rect 457774 278858 457946 279094
rect 458182 278858 458354 279094
rect 457774 243414 458354 278858
rect 457774 243178 457946 243414
rect 458182 243178 458354 243414
rect 457774 243094 458354 243178
rect 457774 242858 457946 243094
rect 458182 242858 458354 243094
rect 457774 207414 458354 242858
rect 457774 207178 457946 207414
rect 458182 207178 458354 207414
rect 457774 207094 458354 207178
rect 457774 206858 457946 207094
rect 458182 206858 458354 207094
rect 457774 171414 458354 206858
rect 457774 171178 457946 171414
rect 458182 171178 458354 171414
rect 457774 171094 458354 171178
rect 457774 170858 457946 171094
rect 458182 170858 458354 171094
rect 457774 135414 458354 170858
rect 457774 135178 457946 135414
rect 458182 135178 458354 135414
rect 457774 135094 458354 135178
rect 457774 134858 457946 135094
rect 458182 134858 458354 135094
rect 457774 99414 458354 134858
rect 457774 99178 457946 99414
rect 458182 99178 458354 99414
rect 457774 99094 458354 99178
rect 457774 98858 457946 99094
rect 458182 98858 458354 99094
rect 457774 63414 458354 98858
rect 457774 63178 457946 63414
rect 458182 63178 458354 63414
rect 457774 63094 458354 63178
rect 457774 62858 457946 63094
rect 458182 62858 458354 63094
rect 457774 27414 458354 62858
rect 457774 27178 457946 27414
rect 458182 27178 458354 27414
rect 457774 27094 458354 27178
rect 457774 26858 457946 27094
rect 458182 26858 458354 27094
rect 457774 -4946 458354 26858
rect 457774 -5182 457946 -4946
rect 458182 -5182 458354 -4946
rect 457774 -5266 458354 -5182
rect 457774 -5502 457946 -5266
rect 458182 -5502 458354 -5266
rect 457774 -5514 458354 -5502
rect 461254 678894 461834 710722
rect 479254 710358 479834 711290
rect 479254 710122 479426 710358
rect 479662 710122 479834 710358
rect 479254 710038 479834 710122
rect 479254 709802 479426 710038
rect 479662 709802 479834 710038
rect 475774 708518 476354 709450
rect 475774 708282 475946 708518
rect 476182 708282 476354 708518
rect 475774 708198 476354 708282
rect 475774 707962 475946 708198
rect 476182 707962 476354 708198
rect 472294 706678 472874 707610
rect 472294 706442 472466 706678
rect 472702 706442 472874 706678
rect 472294 706358 472874 706442
rect 472294 706122 472466 706358
rect 472702 706122 472874 706358
rect 461254 678658 461426 678894
rect 461662 678658 461834 678894
rect 461254 678574 461834 678658
rect 461254 678338 461426 678574
rect 461662 678338 461834 678574
rect 461254 642894 461834 678338
rect 461254 642658 461426 642894
rect 461662 642658 461834 642894
rect 461254 642574 461834 642658
rect 461254 642338 461426 642574
rect 461662 642338 461834 642574
rect 461254 606894 461834 642338
rect 461254 606658 461426 606894
rect 461662 606658 461834 606894
rect 461254 606574 461834 606658
rect 461254 606338 461426 606574
rect 461662 606338 461834 606574
rect 461254 570894 461834 606338
rect 461254 570658 461426 570894
rect 461662 570658 461834 570894
rect 461254 570574 461834 570658
rect 461254 570338 461426 570574
rect 461662 570338 461834 570574
rect 461254 534894 461834 570338
rect 461254 534658 461426 534894
rect 461662 534658 461834 534894
rect 461254 534574 461834 534658
rect 461254 534338 461426 534574
rect 461662 534338 461834 534574
rect 461254 498894 461834 534338
rect 461254 498658 461426 498894
rect 461662 498658 461834 498894
rect 461254 498574 461834 498658
rect 461254 498338 461426 498574
rect 461662 498338 461834 498574
rect 461254 462894 461834 498338
rect 461254 462658 461426 462894
rect 461662 462658 461834 462894
rect 461254 462574 461834 462658
rect 461254 462338 461426 462574
rect 461662 462338 461834 462574
rect 461254 426894 461834 462338
rect 461254 426658 461426 426894
rect 461662 426658 461834 426894
rect 461254 426574 461834 426658
rect 461254 426338 461426 426574
rect 461662 426338 461834 426574
rect 461254 390894 461834 426338
rect 461254 390658 461426 390894
rect 461662 390658 461834 390894
rect 461254 390574 461834 390658
rect 461254 390338 461426 390574
rect 461662 390338 461834 390574
rect 461254 354894 461834 390338
rect 461254 354658 461426 354894
rect 461662 354658 461834 354894
rect 461254 354574 461834 354658
rect 461254 354338 461426 354574
rect 461662 354338 461834 354574
rect 461254 318894 461834 354338
rect 461254 318658 461426 318894
rect 461662 318658 461834 318894
rect 461254 318574 461834 318658
rect 461254 318338 461426 318574
rect 461662 318338 461834 318574
rect 461254 282894 461834 318338
rect 461254 282658 461426 282894
rect 461662 282658 461834 282894
rect 461254 282574 461834 282658
rect 461254 282338 461426 282574
rect 461662 282338 461834 282574
rect 461254 246894 461834 282338
rect 461254 246658 461426 246894
rect 461662 246658 461834 246894
rect 461254 246574 461834 246658
rect 461254 246338 461426 246574
rect 461662 246338 461834 246574
rect 461254 210894 461834 246338
rect 461254 210658 461426 210894
rect 461662 210658 461834 210894
rect 461254 210574 461834 210658
rect 461254 210338 461426 210574
rect 461662 210338 461834 210574
rect 461254 174894 461834 210338
rect 461254 174658 461426 174894
rect 461662 174658 461834 174894
rect 461254 174574 461834 174658
rect 461254 174338 461426 174574
rect 461662 174338 461834 174574
rect 461254 138894 461834 174338
rect 461254 138658 461426 138894
rect 461662 138658 461834 138894
rect 461254 138574 461834 138658
rect 461254 138338 461426 138574
rect 461662 138338 461834 138574
rect 461254 102894 461834 138338
rect 461254 102658 461426 102894
rect 461662 102658 461834 102894
rect 461254 102574 461834 102658
rect 461254 102338 461426 102574
rect 461662 102338 461834 102574
rect 461254 66894 461834 102338
rect 461254 66658 461426 66894
rect 461662 66658 461834 66894
rect 461254 66574 461834 66658
rect 461254 66338 461426 66574
rect 461662 66338 461834 66574
rect 461254 30894 461834 66338
rect 461254 30658 461426 30894
rect 461662 30658 461834 30894
rect 461254 30574 461834 30658
rect 461254 30338 461426 30574
rect 461662 30338 461834 30574
rect 443254 -6102 443426 -5866
rect 443662 -6102 443834 -5866
rect 443254 -6186 443834 -6102
rect 443254 -6422 443426 -6186
rect 443662 -6422 443834 -6186
rect 443254 -7354 443834 -6422
rect 461254 -6786 461834 30338
rect 468814 704838 469394 705770
rect 468814 704602 468986 704838
rect 469222 704602 469394 704838
rect 468814 704518 469394 704602
rect 468814 704282 468986 704518
rect 469222 704282 469394 704518
rect 468814 686454 469394 704282
rect 468814 686218 468986 686454
rect 469222 686218 469394 686454
rect 468814 686134 469394 686218
rect 468814 685898 468986 686134
rect 469222 685898 469394 686134
rect 468814 650454 469394 685898
rect 468814 650218 468986 650454
rect 469222 650218 469394 650454
rect 468814 650134 469394 650218
rect 468814 649898 468986 650134
rect 469222 649898 469394 650134
rect 468814 614454 469394 649898
rect 468814 614218 468986 614454
rect 469222 614218 469394 614454
rect 468814 614134 469394 614218
rect 468814 613898 468986 614134
rect 469222 613898 469394 614134
rect 468814 578454 469394 613898
rect 468814 578218 468986 578454
rect 469222 578218 469394 578454
rect 468814 578134 469394 578218
rect 468814 577898 468986 578134
rect 469222 577898 469394 578134
rect 468814 542454 469394 577898
rect 468814 542218 468986 542454
rect 469222 542218 469394 542454
rect 468814 542134 469394 542218
rect 468814 541898 468986 542134
rect 469222 541898 469394 542134
rect 468814 506454 469394 541898
rect 468814 506218 468986 506454
rect 469222 506218 469394 506454
rect 468814 506134 469394 506218
rect 468814 505898 468986 506134
rect 469222 505898 469394 506134
rect 468814 470454 469394 505898
rect 468814 470218 468986 470454
rect 469222 470218 469394 470454
rect 468814 470134 469394 470218
rect 468814 469898 468986 470134
rect 469222 469898 469394 470134
rect 468814 434454 469394 469898
rect 468814 434218 468986 434454
rect 469222 434218 469394 434454
rect 468814 434134 469394 434218
rect 468814 433898 468986 434134
rect 469222 433898 469394 434134
rect 468814 398454 469394 433898
rect 468814 398218 468986 398454
rect 469222 398218 469394 398454
rect 468814 398134 469394 398218
rect 468814 397898 468986 398134
rect 469222 397898 469394 398134
rect 468814 362454 469394 397898
rect 468814 362218 468986 362454
rect 469222 362218 469394 362454
rect 468814 362134 469394 362218
rect 468814 361898 468986 362134
rect 469222 361898 469394 362134
rect 468814 326454 469394 361898
rect 468814 326218 468986 326454
rect 469222 326218 469394 326454
rect 468814 326134 469394 326218
rect 468814 325898 468986 326134
rect 469222 325898 469394 326134
rect 468814 290454 469394 325898
rect 468814 290218 468986 290454
rect 469222 290218 469394 290454
rect 468814 290134 469394 290218
rect 468814 289898 468986 290134
rect 469222 289898 469394 290134
rect 468814 254454 469394 289898
rect 468814 254218 468986 254454
rect 469222 254218 469394 254454
rect 468814 254134 469394 254218
rect 468814 253898 468986 254134
rect 469222 253898 469394 254134
rect 468814 218454 469394 253898
rect 468814 218218 468986 218454
rect 469222 218218 469394 218454
rect 468814 218134 469394 218218
rect 468814 217898 468986 218134
rect 469222 217898 469394 218134
rect 468814 182454 469394 217898
rect 468814 182218 468986 182454
rect 469222 182218 469394 182454
rect 468814 182134 469394 182218
rect 468814 181898 468986 182134
rect 469222 181898 469394 182134
rect 468814 146454 469394 181898
rect 468814 146218 468986 146454
rect 469222 146218 469394 146454
rect 468814 146134 469394 146218
rect 468814 145898 468986 146134
rect 469222 145898 469394 146134
rect 468814 110454 469394 145898
rect 468814 110218 468986 110454
rect 469222 110218 469394 110454
rect 468814 110134 469394 110218
rect 468814 109898 468986 110134
rect 469222 109898 469394 110134
rect 468814 74454 469394 109898
rect 468814 74218 468986 74454
rect 469222 74218 469394 74454
rect 468814 74134 469394 74218
rect 468814 73898 468986 74134
rect 469222 73898 469394 74134
rect 468814 38454 469394 73898
rect 468814 38218 468986 38454
rect 469222 38218 469394 38454
rect 468814 38134 469394 38218
rect 468814 37898 468986 38134
rect 469222 37898 469394 38134
rect 468814 2454 469394 37898
rect 468814 2218 468986 2454
rect 469222 2218 469394 2454
rect 468814 2134 469394 2218
rect 468814 1898 468986 2134
rect 469222 1898 469394 2134
rect 468814 -346 469394 1898
rect 468814 -582 468986 -346
rect 469222 -582 469394 -346
rect 468814 -666 469394 -582
rect 468814 -902 468986 -666
rect 469222 -902 469394 -666
rect 468814 -1834 469394 -902
rect 472294 689934 472874 706122
rect 472294 689698 472466 689934
rect 472702 689698 472874 689934
rect 472294 689614 472874 689698
rect 472294 689378 472466 689614
rect 472702 689378 472874 689614
rect 472294 653934 472874 689378
rect 472294 653698 472466 653934
rect 472702 653698 472874 653934
rect 472294 653614 472874 653698
rect 472294 653378 472466 653614
rect 472702 653378 472874 653614
rect 472294 617934 472874 653378
rect 472294 617698 472466 617934
rect 472702 617698 472874 617934
rect 472294 617614 472874 617698
rect 472294 617378 472466 617614
rect 472702 617378 472874 617614
rect 472294 581934 472874 617378
rect 472294 581698 472466 581934
rect 472702 581698 472874 581934
rect 472294 581614 472874 581698
rect 472294 581378 472466 581614
rect 472702 581378 472874 581614
rect 472294 545934 472874 581378
rect 472294 545698 472466 545934
rect 472702 545698 472874 545934
rect 472294 545614 472874 545698
rect 472294 545378 472466 545614
rect 472702 545378 472874 545614
rect 472294 509934 472874 545378
rect 472294 509698 472466 509934
rect 472702 509698 472874 509934
rect 472294 509614 472874 509698
rect 472294 509378 472466 509614
rect 472702 509378 472874 509614
rect 472294 473934 472874 509378
rect 472294 473698 472466 473934
rect 472702 473698 472874 473934
rect 472294 473614 472874 473698
rect 472294 473378 472466 473614
rect 472702 473378 472874 473614
rect 472294 437934 472874 473378
rect 472294 437698 472466 437934
rect 472702 437698 472874 437934
rect 472294 437614 472874 437698
rect 472294 437378 472466 437614
rect 472702 437378 472874 437614
rect 472294 401934 472874 437378
rect 472294 401698 472466 401934
rect 472702 401698 472874 401934
rect 472294 401614 472874 401698
rect 472294 401378 472466 401614
rect 472702 401378 472874 401614
rect 472294 365934 472874 401378
rect 472294 365698 472466 365934
rect 472702 365698 472874 365934
rect 472294 365614 472874 365698
rect 472294 365378 472466 365614
rect 472702 365378 472874 365614
rect 472294 329934 472874 365378
rect 472294 329698 472466 329934
rect 472702 329698 472874 329934
rect 472294 329614 472874 329698
rect 472294 329378 472466 329614
rect 472702 329378 472874 329614
rect 472294 293934 472874 329378
rect 472294 293698 472466 293934
rect 472702 293698 472874 293934
rect 472294 293614 472874 293698
rect 472294 293378 472466 293614
rect 472702 293378 472874 293614
rect 472294 257934 472874 293378
rect 472294 257698 472466 257934
rect 472702 257698 472874 257934
rect 472294 257614 472874 257698
rect 472294 257378 472466 257614
rect 472702 257378 472874 257614
rect 472294 221934 472874 257378
rect 472294 221698 472466 221934
rect 472702 221698 472874 221934
rect 472294 221614 472874 221698
rect 472294 221378 472466 221614
rect 472702 221378 472874 221614
rect 472294 185934 472874 221378
rect 472294 185698 472466 185934
rect 472702 185698 472874 185934
rect 472294 185614 472874 185698
rect 472294 185378 472466 185614
rect 472702 185378 472874 185614
rect 472294 149934 472874 185378
rect 472294 149698 472466 149934
rect 472702 149698 472874 149934
rect 472294 149614 472874 149698
rect 472294 149378 472466 149614
rect 472702 149378 472874 149614
rect 472294 113934 472874 149378
rect 472294 113698 472466 113934
rect 472702 113698 472874 113934
rect 472294 113614 472874 113698
rect 472294 113378 472466 113614
rect 472702 113378 472874 113614
rect 472294 77934 472874 113378
rect 472294 77698 472466 77934
rect 472702 77698 472874 77934
rect 472294 77614 472874 77698
rect 472294 77378 472466 77614
rect 472702 77378 472874 77614
rect 472294 41934 472874 77378
rect 472294 41698 472466 41934
rect 472702 41698 472874 41934
rect 472294 41614 472874 41698
rect 472294 41378 472466 41614
rect 472702 41378 472874 41614
rect 472294 5934 472874 41378
rect 472294 5698 472466 5934
rect 472702 5698 472874 5934
rect 472294 5614 472874 5698
rect 472294 5378 472466 5614
rect 472702 5378 472874 5614
rect 472294 -2186 472874 5378
rect 472294 -2422 472466 -2186
rect 472702 -2422 472874 -2186
rect 472294 -2506 472874 -2422
rect 472294 -2742 472466 -2506
rect 472702 -2742 472874 -2506
rect 472294 -3674 472874 -2742
rect 475774 693414 476354 707962
rect 475774 693178 475946 693414
rect 476182 693178 476354 693414
rect 475774 693094 476354 693178
rect 475774 692858 475946 693094
rect 476182 692858 476354 693094
rect 475774 657414 476354 692858
rect 475774 657178 475946 657414
rect 476182 657178 476354 657414
rect 475774 657094 476354 657178
rect 475774 656858 475946 657094
rect 476182 656858 476354 657094
rect 475774 621414 476354 656858
rect 475774 621178 475946 621414
rect 476182 621178 476354 621414
rect 475774 621094 476354 621178
rect 475774 620858 475946 621094
rect 476182 620858 476354 621094
rect 475774 585414 476354 620858
rect 475774 585178 475946 585414
rect 476182 585178 476354 585414
rect 475774 585094 476354 585178
rect 475774 584858 475946 585094
rect 476182 584858 476354 585094
rect 475774 549414 476354 584858
rect 475774 549178 475946 549414
rect 476182 549178 476354 549414
rect 475774 549094 476354 549178
rect 475774 548858 475946 549094
rect 476182 548858 476354 549094
rect 475774 513414 476354 548858
rect 475774 513178 475946 513414
rect 476182 513178 476354 513414
rect 475774 513094 476354 513178
rect 475774 512858 475946 513094
rect 476182 512858 476354 513094
rect 475774 477414 476354 512858
rect 475774 477178 475946 477414
rect 476182 477178 476354 477414
rect 475774 477094 476354 477178
rect 475774 476858 475946 477094
rect 476182 476858 476354 477094
rect 475774 441414 476354 476858
rect 475774 441178 475946 441414
rect 476182 441178 476354 441414
rect 475774 441094 476354 441178
rect 475774 440858 475946 441094
rect 476182 440858 476354 441094
rect 475774 405414 476354 440858
rect 475774 405178 475946 405414
rect 476182 405178 476354 405414
rect 475774 405094 476354 405178
rect 475774 404858 475946 405094
rect 476182 404858 476354 405094
rect 475774 369414 476354 404858
rect 475774 369178 475946 369414
rect 476182 369178 476354 369414
rect 475774 369094 476354 369178
rect 475774 368858 475946 369094
rect 476182 368858 476354 369094
rect 475774 333414 476354 368858
rect 475774 333178 475946 333414
rect 476182 333178 476354 333414
rect 475774 333094 476354 333178
rect 475774 332858 475946 333094
rect 476182 332858 476354 333094
rect 475774 297414 476354 332858
rect 475774 297178 475946 297414
rect 476182 297178 476354 297414
rect 475774 297094 476354 297178
rect 475774 296858 475946 297094
rect 476182 296858 476354 297094
rect 475774 261414 476354 296858
rect 475774 261178 475946 261414
rect 476182 261178 476354 261414
rect 475774 261094 476354 261178
rect 475774 260858 475946 261094
rect 476182 260858 476354 261094
rect 475774 225414 476354 260858
rect 475774 225178 475946 225414
rect 476182 225178 476354 225414
rect 475774 225094 476354 225178
rect 475774 224858 475946 225094
rect 476182 224858 476354 225094
rect 475774 189414 476354 224858
rect 475774 189178 475946 189414
rect 476182 189178 476354 189414
rect 475774 189094 476354 189178
rect 475774 188858 475946 189094
rect 476182 188858 476354 189094
rect 475774 153414 476354 188858
rect 475774 153178 475946 153414
rect 476182 153178 476354 153414
rect 475774 153094 476354 153178
rect 475774 152858 475946 153094
rect 476182 152858 476354 153094
rect 475774 117414 476354 152858
rect 475774 117178 475946 117414
rect 476182 117178 476354 117414
rect 475774 117094 476354 117178
rect 475774 116858 475946 117094
rect 476182 116858 476354 117094
rect 475774 81414 476354 116858
rect 475774 81178 475946 81414
rect 476182 81178 476354 81414
rect 475774 81094 476354 81178
rect 475774 80858 475946 81094
rect 476182 80858 476354 81094
rect 475774 45414 476354 80858
rect 475774 45178 475946 45414
rect 476182 45178 476354 45414
rect 475774 45094 476354 45178
rect 475774 44858 475946 45094
rect 476182 44858 476354 45094
rect 475774 9414 476354 44858
rect 475774 9178 475946 9414
rect 476182 9178 476354 9414
rect 475774 9094 476354 9178
rect 475774 8858 475946 9094
rect 476182 8858 476354 9094
rect 475774 -4026 476354 8858
rect 475774 -4262 475946 -4026
rect 476182 -4262 476354 -4026
rect 475774 -4346 476354 -4262
rect 475774 -4582 475946 -4346
rect 476182 -4582 476354 -4346
rect 475774 -5514 476354 -4582
rect 479254 696894 479834 709802
rect 497254 711278 497834 711290
rect 497254 711042 497426 711278
rect 497662 711042 497834 711278
rect 497254 710958 497834 711042
rect 497254 710722 497426 710958
rect 497662 710722 497834 710958
rect 493774 709438 494354 709450
rect 493774 709202 493946 709438
rect 494182 709202 494354 709438
rect 493774 709118 494354 709202
rect 493774 708882 493946 709118
rect 494182 708882 494354 709118
rect 490294 707598 490874 707610
rect 490294 707362 490466 707598
rect 490702 707362 490874 707598
rect 490294 707278 490874 707362
rect 490294 707042 490466 707278
rect 490702 707042 490874 707278
rect 479254 696658 479426 696894
rect 479662 696658 479834 696894
rect 479254 696574 479834 696658
rect 479254 696338 479426 696574
rect 479662 696338 479834 696574
rect 479254 660894 479834 696338
rect 479254 660658 479426 660894
rect 479662 660658 479834 660894
rect 479254 660574 479834 660658
rect 479254 660338 479426 660574
rect 479662 660338 479834 660574
rect 479254 624894 479834 660338
rect 479254 624658 479426 624894
rect 479662 624658 479834 624894
rect 479254 624574 479834 624658
rect 479254 624338 479426 624574
rect 479662 624338 479834 624574
rect 479254 588894 479834 624338
rect 479254 588658 479426 588894
rect 479662 588658 479834 588894
rect 479254 588574 479834 588658
rect 479254 588338 479426 588574
rect 479662 588338 479834 588574
rect 479254 552894 479834 588338
rect 479254 552658 479426 552894
rect 479662 552658 479834 552894
rect 479254 552574 479834 552658
rect 479254 552338 479426 552574
rect 479662 552338 479834 552574
rect 479254 516894 479834 552338
rect 479254 516658 479426 516894
rect 479662 516658 479834 516894
rect 479254 516574 479834 516658
rect 479254 516338 479426 516574
rect 479662 516338 479834 516574
rect 479254 480894 479834 516338
rect 479254 480658 479426 480894
rect 479662 480658 479834 480894
rect 479254 480574 479834 480658
rect 479254 480338 479426 480574
rect 479662 480338 479834 480574
rect 479254 444894 479834 480338
rect 479254 444658 479426 444894
rect 479662 444658 479834 444894
rect 479254 444574 479834 444658
rect 479254 444338 479426 444574
rect 479662 444338 479834 444574
rect 479254 408894 479834 444338
rect 479254 408658 479426 408894
rect 479662 408658 479834 408894
rect 479254 408574 479834 408658
rect 479254 408338 479426 408574
rect 479662 408338 479834 408574
rect 479254 372894 479834 408338
rect 479254 372658 479426 372894
rect 479662 372658 479834 372894
rect 479254 372574 479834 372658
rect 479254 372338 479426 372574
rect 479662 372338 479834 372574
rect 479254 336894 479834 372338
rect 479254 336658 479426 336894
rect 479662 336658 479834 336894
rect 479254 336574 479834 336658
rect 479254 336338 479426 336574
rect 479662 336338 479834 336574
rect 479254 300894 479834 336338
rect 479254 300658 479426 300894
rect 479662 300658 479834 300894
rect 479254 300574 479834 300658
rect 479254 300338 479426 300574
rect 479662 300338 479834 300574
rect 479254 264894 479834 300338
rect 479254 264658 479426 264894
rect 479662 264658 479834 264894
rect 479254 264574 479834 264658
rect 479254 264338 479426 264574
rect 479662 264338 479834 264574
rect 479254 228894 479834 264338
rect 479254 228658 479426 228894
rect 479662 228658 479834 228894
rect 479254 228574 479834 228658
rect 479254 228338 479426 228574
rect 479662 228338 479834 228574
rect 479254 192894 479834 228338
rect 479254 192658 479426 192894
rect 479662 192658 479834 192894
rect 479254 192574 479834 192658
rect 479254 192338 479426 192574
rect 479662 192338 479834 192574
rect 479254 156894 479834 192338
rect 479254 156658 479426 156894
rect 479662 156658 479834 156894
rect 479254 156574 479834 156658
rect 479254 156338 479426 156574
rect 479662 156338 479834 156574
rect 479254 120894 479834 156338
rect 479254 120658 479426 120894
rect 479662 120658 479834 120894
rect 479254 120574 479834 120658
rect 479254 120338 479426 120574
rect 479662 120338 479834 120574
rect 479254 84894 479834 120338
rect 479254 84658 479426 84894
rect 479662 84658 479834 84894
rect 479254 84574 479834 84658
rect 479254 84338 479426 84574
rect 479662 84338 479834 84574
rect 479254 48894 479834 84338
rect 479254 48658 479426 48894
rect 479662 48658 479834 48894
rect 479254 48574 479834 48658
rect 479254 48338 479426 48574
rect 479662 48338 479834 48574
rect 479254 12894 479834 48338
rect 479254 12658 479426 12894
rect 479662 12658 479834 12894
rect 479254 12574 479834 12658
rect 479254 12338 479426 12574
rect 479662 12338 479834 12574
rect 461254 -7022 461426 -6786
rect 461662 -7022 461834 -6786
rect 461254 -7106 461834 -7022
rect 461254 -7342 461426 -7106
rect 461662 -7342 461834 -7106
rect 461254 -7354 461834 -7342
rect 479254 -5866 479834 12338
rect 486814 705758 487394 705770
rect 486814 705522 486986 705758
rect 487222 705522 487394 705758
rect 486814 705438 487394 705522
rect 486814 705202 486986 705438
rect 487222 705202 487394 705438
rect 486814 668454 487394 705202
rect 486814 668218 486986 668454
rect 487222 668218 487394 668454
rect 486814 668134 487394 668218
rect 486814 667898 486986 668134
rect 487222 667898 487394 668134
rect 486814 632454 487394 667898
rect 486814 632218 486986 632454
rect 487222 632218 487394 632454
rect 486814 632134 487394 632218
rect 486814 631898 486986 632134
rect 487222 631898 487394 632134
rect 486814 596454 487394 631898
rect 486814 596218 486986 596454
rect 487222 596218 487394 596454
rect 486814 596134 487394 596218
rect 486814 595898 486986 596134
rect 487222 595898 487394 596134
rect 486814 560454 487394 595898
rect 486814 560218 486986 560454
rect 487222 560218 487394 560454
rect 486814 560134 487394 560218
rect 486814 559898 486986 560134
rect 487222 559898 487394 560134
rect 486814 524454 487394 559898
rect 486814 524218 486986 524454
rect 487222 524218 487394 524454
rect 486814 524134 487394 524218
rect 486814 523898 486986 524134
rect 487222 523898 487394 524134
rect 486814 488454 487394 523898
rect 486814 488218 486986 488454
rect 487222 488218 487394 488454
rect 486814 488134 487394 488218
rect 486814 487898 486986 488134
rect 487222 487898 487394 488134
rect 486814 452454 487394 487898
rect 486814 452218 486986 452454
rect 487222 452218 487394 452454
rect 486814 452134 487394 452218
rect 486814 451898 486986 452134
rect 487222 451898 487394 452134
rect 486814 416454 487394 451898
rect 486814 416218 486986 416454
rect 487222 416218 487394 416454
rect 486814 416134 487394 416218
rect 486814 415898 486986 416134
rect 487222 415898 487394 416134
rect 486814 380454 487394 415898
rect 486814 380218 486986 380454
rect 487222 380218 487394 380454
rect 486814 380134 487394 380218
rect 486814 379898 486986 380134
rect 487222 379898 487394 380134
rect 486814 344454 487394 379898
rect 486814 344218 486986 344454
rect 487222 344218 487394 344454
rect 486814 344134 487394 344218
rect 486814 343898 486986 344134
rect 487222 343898 487394 344134
rect 486814 308454 487394 343898
rect 486814 308218 486986 308454
rect 487222 308218 487394 308454
rect 486814 308134 487394 308218
rect 486814 307898 486986 308134
rect 487222 307898 487394 308134
rect 486814 272454 487394 307898
rect 486814 272218 486986 272454
rect 487222 272218 487394 272454
rect 486814 272134 487394 272218
rect 486814 271898 486986 272134
rect 487222 271898 487394 272134
rect 486814 236454 487394 271898
rect 486814 236218 486986 236454
rect 487222 236218 487394 236454
rect 486814 236134 487394 236218
rect 486814 235898 486986 236134
rect 487222 235898 487394 236134
rect 486814 200454 487394 235898
rect 486814 200218 486986 200454
rect 487222 200218 487394 200454
rect 486814 200134 487394 200218
rect 486814 199898 486986 200134
rect 487222 199898 487394 200134
rect 486814 164454 487394 199898
rect 486814 164218 486986 164454
rect 487222 164218 487394 164454
rect 486814 164134 487394 164218
rect 486814 163898 486986 164134
rect 487222 163898 487394 164134
rect 486814 128454 487394 163898
rect 486814 128218 486986 128454
rect 487222 128218 487394 128454
rect 486814 128134 487394 128218
rect 486814 127898 486986 128134
rect 487222 127898 487394 128134
rect 486814 92454 487394 127898
rect 486814 92218 486986 92454
rect 487222 92218 487394 92454
rect 486814 92134 487394 92218
rect 486814 91898 486986 92134
rect 487222 91898 487394 92134
rect 486814 56454 487394 91898
rect 486814 56218 486986 56454
rect 487222 56218 487394 56454
rect 486814 56134 487394 56218
rect 486814 55898 486986 56134
rect 487222 55898 487394 56134
rect 486814 20454 487394 55898
rect 486814 20218 486986 20454
rect 487222 20218 487394 20454
rect 486814 20134 487394 20218
rect 486814 19898 486986 20134
rect 487222 19898 487394 20134
rect 486814 -1266 487394 19898
rect 486814 -1502 486986 -1266
rect 487222 -1502 487394 -1266
rect 486814 -1586 487394 -1502
rect 486814 -1822 486986 -1586
rect 487222 -1822 487394 -1586
rect 486814 -1834 487394 -1822
rect 490294 671934 490874 707042
rect 490294 671698 490466 671934
rect 490702 671698 490874 671934
rect 490294 671614 490874 671698
rect 490294 671378 490466 671614
rect 490702 671378 490874 671614
rect 490294 635934 490874 671378
rect 490294 635698 490466 635934
rect 490702 635698 490874 635934
rect 490294 635614 490874 635698
rect 490294 635378 490466 635614
rect 490702 635378 490874 635614
rect 490294 599934 490874 635378
rect 490294 599698 490466 599934
rect 490702 599698 490874 599934
rect 490294 599614 490874 599698
rect 490294 599378 490466 599614
rect 490702 599378 490874 599614
rect 490294 563934 490874 599378
rect 490294 563698 490466 563934
rect 490702 563698 490874 563934
rect 490294 563614 490874 563698
rect 490294 563378 490466 563614
rect 490702 563378 490874 563614
rect 490294 527934 490874 563378
rect 490294 527698 490466 527934
rect 490702 527698 490874 527934
rect 490294 527614 490874 527698
rect 490294 527378 490466 527614
rect 490702 527378 490874 527614
rect 490294 491934 490874 527378
rect 490294 491698 490466 491934
rect 490702 491698 490874 491934
rect 490294 491614 490874 491698
rect 490294 491378 490466 491614
rect 490702 491378 490874 491614
rect 490294 455934 490874 491378
rect 490294 455698 490466 455934
rect 490702 455698 490874 455934
rect 490294 455614 490874 455698
rect 490294 455378 490466 455614
rect 490702 455378 490874 455614
rect 490294 419934 490874 455378
rect 490294 419698 490466 419934
rect 490702 419698 490874 419934
rect 490294 419614 490874 419698
rect 490294 419378 490466 419614
rect 490702 419378 490874 419614
rect 490294 383934 490874 419378
rect 490294 383698 490466 383934
rect 490702 383698 490874 383934
rect 490294 383614 490874 383698
rect 490294 383378 490466 383614
rect 490702 383378 490874 383614
rect 490294 347934 490874 383378
rect 490294 347698 490466 347934
rect 490702 347698 490874 347934
rect 490294 347614 490874 347698
rect 490294 347378 490466 347614
rect 490702 347378 490874 347614
rect 490294 311934 490874 347378
rect 490294 311698 490466 311934
rect 490702 311698 490874 311934
rect 490294 311614 490874 311698
rect 490294 311378 490466 311614
rect 490702 311378 490874 311614
rect 490294 275934 490874 311378
rect 490294 275698 490466 275934
rect 490702 275698 490874 275934
rect 490294 275614 490874 275698
rect 490294 275378 490466 275614
rect 490702 275378 490874 275614
rect 490294 239934 490874 275378
rect 490294 239698 490466 239934
rect 490702 239698 490874 239934
rect 490294 239614 490874 239698
rect 490294 239378 490466 239614
rect 490702 239378 490874 239614
rect 490294 203934 490874 239378
rect 490294 203698 490466 203934
rect 490702 203698 490874 203934
rect 490294 203614 490874 203698
rect 490294 203378 490466 203614
rect 490702 203378 490874 203614
rect 490294 167934 490874 203378
rect 490294 167698 490466 167934
rect 490702 167698 490874 167934
rect 490294 167614 490874 167698
rect 490294 167378 490466 167614
rect 490702 167378 490874 167614
rect 490294 131934 490874 167378
rect 490294 131698 490466 131934
rect 490702 131698 490874 131934
rect 490294 131614 490874 131698
rect 490294 131378 490466 131614
rect 490702 131378 490874 131614
rect 490294 95934 490874 131378
rect 490294 95698 490466 95934
rect 490702 95698 490874 95934
rect 490294 95614 490874 95698
rect 490294 95378 490466 95614
rect 490702 95378 490874 95614
rect 490294 59934 490874 95378
rect 490294 59698 490466 59934
rect 490702 59698 490874 59934
rect 490294 59614 490874 59698
rect 490294 59378 490466 59614
rect 490702 59378 490874 59614
rect 490294 23934 490874 59378
rect 490294 23698 490466 23934
rect 490702 23698 490874 23934
rect 490294 23614 490874 23698
rect 490294 23378 490466 23614
rect 490702 23378 490874 23614
rect 490294 -3106 490874 23378
rect 490294 -3342 490466 -3106
rect 490702 -3342 490874 -3106
rect 490294 -3426 490874 -3342
rect 490294 -3662 490466 -3426
rect 490702 -3662 490874 -3426
rect 490294 -3674 490874 -3662
rect 493774 675414 494354 708882
rect 493774 675178 493946 675414
rect 494182 675178 494354 675414
rect 493774 675094 494354 675178
rect 493774 674858 493946 675094
rect 494182 674858 494354 675094
rect 493774 639414 494354 674858
rect 493774 639178 493946 639414
rect 494182 639178 494354 639414
rect 493774 639094 494354 639178
rect 493774 638858 493946 639094
rect 494182 638858 494354 639094
rect 493774 603414 494354 638858
rect 493774 603178 493946 603414
rect 494182 603178 494354 603414
rect 493774 603094 494354 603178
rect 493774 602858 493946 603094
rect 494182 602858 494354 603094
rect 493774 567414 494354 602858
rect 493774 567178 493946 567414
rect 494182 567178 494354 567414
rect 493774 567094 494354 567178
rect 493774 566858 493946 567094
rect 494182 566858 494354 567094
rect 493774 531414 494354 566858
rect 493774 531178 493946 531414
rect 494182 531178 494354 531414
rect 493774 531094 494354 531178
rect 493774 530858 493946 531094
rect 494182 530858 494354 531094
rect 493774 495414 494354 530858
rect 493774 495178 493946 495414
rect 494182 495178 494354 495414
rect 493774 495094 494354 495178
rect 493774 494858 493946 495094
rect 494182 494858 494354 495094
rect 493774 459414 494354 494858
rect 493774 459178 493946 459414
rect 494182 459178 494354 459414
rect 493774 459094 494354 459178
rect 493774 458858 493946 459094
rect 494182 458858 494354 459094
rect 493774 423414 494354 458858
rect 493774 423178 493946 423414
rect 494182 423178 494354 423414
rect 493774 423094 494354 423178
rect 493774 422858 493946 423094
rect 494182 422858 494354 423094
rect 493774 387414 494354 422858
rect 493774 387178 493946 387414
rect 494182 387178 494354 387414
rect 493774 387094 494354 387178
rect 493774 386858 493946 387094
rect 494182 386858 494354 387094
rect 493774 351414 494354 386858
rect 493774 351178 493946 351414
rect 494182 351178 494354 351414
rect 493774 351094 494354 351178
rect 493774 350858 493946 351094
rect 494182 350858 494354 351094
rect 493774 315414 494354 350858
rect 493774 315178 493946 315414
rect 494182 315178 494354 315414
rect 493774 315094 494354 315178
rect 493774 314858 493946 315094
rect 494182 314858 494354 315094
rect 493774 279414 494354 314858
rect 493774 279178 493946 279414
rect 494182 279178 494354 279414
rect 493774 279094 494354 279178
rect 493774 278858 493946 279094
rect 494182 278858 494354 279094
rect 493774 243414 494354 278858
rect 493774 243178 493946 243414
rect 494182 243178 494354 243414
rect 493774 243094 494354 243178
rect 493774 242858 493946 243094
rect 494182 242858 494354 243094
rect 493774 207414 494354 242858
rect 493774 207178 493946 207414
rect 494182 207178 494354 207414
rect 493774 207094 494354 207178
rect 493774 206858 493946 207094
rect 494182 206858 494354 207094
rect 493774 171414 494354 206858
rect 493774 171178 493946 171414
rect 494182 171178 494354 171414
rect 493774 171094 494354 171178
rect 493774 170858 493946 171094
rect 494182 170858 494354 171094
rect 493774 135414 494354 170858
rect 493774 135178 493946 135414
rect 494182 135178 494354 135414
rect 493774 135094 494354 135178
rect 493774 134858 493946 135094
rect 494182 134858 494354 135094
rect 493774 99414 494354 134858
rect 493774 99178 493946 99414
rect 494182 99178 494354 99414
rect 493774 99094 494354 99178
rect 493774 98858 493946 99094
rect 494182 98858 494354 99094
rect 493774 63414 494354 98858
rect 493774 63178 493946 63414
rect 494182 63178 494354 63414
rect 493774 63094 494354 63178
rect 493774 62858 493946 63094
rect 494182 62858 494354 63094
rect 493774 27414 494354 62858
rect 493774 27178 493946 27414
rect 494182 27178 494354 27414
rect 493774 27094 494354 27178
rect 493774 26858 493946 27094
rect 494182 26858 494354 27094
rect 493774 -4946 494354 26858
rect 493774 -5182 493946 -4946
rect 494182 -5182 494354 -4946
rect 493774 -5266 494354 -5182
rect 493774 -5502 493946 -5266
rect 494182 -5502 494354 -5266
rect 493774 -5514 494354 -5502
rect 497254 678894 497834 710722
rect 515254 710358 515834 711290
rect 515254 710122 515426 710358
rect 515662 710122 515834 710358
rect 515254 710038 515834 710122
rect 515254 709802 515426 710038
rect 515662 709802 515834 710038
rect 511774 708518 512354 709450
rect 511774 708282 511946 708518
rect 512182 708282 512354 708518
rect 511774 708198 512354 708282
rect 511774 707962 511946 708198
rect 512182 707962 512354 708198
rect 508294 706678 508874 707610
rect 508294 706442 508466 706678
rect 508702 706442 508874 706678
rect 508294 706358 508874 706442
rect 508294 706122 508466 706358
rect 508702 706122 508874 706358
rect 497254 678658 497426 678894
rect 497662 678658 497834 678894
rect 497254 678574 497834 678658
rect 497254 678338 497426 678574
rect 497662 678338 497834 678574
rect 497254 642894 497834 678338
rect 497254 642658 497426 642894
rect 497662 642658 497834 642894
rect 497254 642574 497834 642658
rect 497254 642338 497426 642574
rect 497662 642338 497834 642574
rect 497254 606894 497834 642338
rect 497254 606658 497426 606894
rect 497662 606658 497834 606894
rect 497254 606574 497834 606658
rect 497254 606338 497426 606574
rect 497662 606338 497834 606574
rect 497254 570894 497834 606338
rect 497254 570658 497426 570894
rect 497662 570658 497834 570894
rect 497254 570574 497834 570658
rect 497254 570338 497426 570574
rect 497662 570338 497834 570574
rect 497254 534894 497834 570338
rect 497254 534658 497426 534894
rect 497662 534658 497834 534894
rect 497254 534574 497834 534658
rect 497254 534338 497426 534574
rect 497662 534338 497834 534574
rect 497254 498894 497834 534338
rect 497254 498658 497426 498894
rect 497662 498658 497834 498894
rect 497254 498574 497834 498658
rect 497254 498338 497426 498574
rect 497662 498338 497834 498574
rect 497254 462894 497834 498338
rect 497254 462658 497426 462894
rect 497662 462658 497834 462894
rect 497254 462574 497834 462658
rect 497254 462338 497426 462574
rect 497662 462338 497834 462574
rect 497254 426894 497834 462338
rect 497254 426658 497426 426894
rect 497662 426658 497834 426894
rect 497254 426574 497834 426658
rect 497254 426338 497426 426574
rect 497662 426338 497834 426574
rect 497254 390894 497834 426338
rect 497254 390658 497426 390894
rect 497662 390658 497834 390894
rect 497254 390574 497834 390658
rect 497254 390338 497426 390574
rect 497662 390338 497834 390574
rect 497254 354894 497834 390338
rect 497254 354658 497426 354894
rect 497662 354658 497834 354894
rect 497254 354574 497834 354658
rect 497254 354338 497426 354574
rect 497662 354338 497834 354574
rect 497254 318894 497834 354338
rect 497254 318658 497426 318894
rect 497662 318658 497834 318894
rect 497254 318574 497834 318658
rect 497254 318338 497426 318574
rect 497662 318338 497834 318574
rect 497254 282894 497834 318338
rect 497254 282658 497426 282894
rect 497662 282658 497834 282894
rect 497254 282574 497834 282658
rect 497254 282338 497426 282574
rect 497662 282338 497834 282574
rect 497254 246894 497834 282338
rect 497254 246658 497426 246894
rect 497662 246658 497834 246894
rect 497254 246574 497834 246658
rect 497254 246338 497426 246574
rect 497662 246338 497834 246574
rect 497254 210894 497834 246338
rect 497254 210658 497426 210894
rect 497662 210658 497834 210894
rect 497254 210574 497834 210658
rect 497254 210338 497426 210574
rect 497662 210338 497834 210574
rect 497254 174894 497834 210338
rect 497254 174658 497426 174894
rect 497662 174658 497834 174894
rect 497254 174574 497834 174658
rect 497254 174338 497426 174574
rect 497662 174338 497834 174574
rect 497254 138894 497834 174338
rect 497254 138658 497426 138894
rect 497662 138658 497834 138894
rect 497254 138574 497834 138658
rect 497254 138338 497426 138574
rect 497662 138338 497834 138574
rect 497254 102894 497834 138338
rect 497254 102658 497426 102894
rect 497662 102658 497834 102894
rect 497254 102574 497834 102658
rect 497254 102338 497426 102574
rect 497662 102338 497834 102574
rect 497254 66894 497834 102338
rect 497254 66658 497426 66894
rect 497662 66658 497834 66894
rect 497254 66574 497834 66658
rect 497254 66338 497426 66574
rect 497662 66338 497834 66574
rect 497254 30894 497834 66338
rect 497254 30658 497426 30894
rect 497662 30658 497834 30894
rect 497254 30574 497834 30658
rect 497254 30338 497426 30574
rect 497662 30338 497834 30574
rect 479254 -6102 479426 -5866
rect 479662 -6102 479834 -5866
rect 479254 -6186 479834 -6102
rect 479254 -6422 479426 -6186
rect 479662 -6422 479834 -6186
rect 479254 -7354 479834 -6422
rect 497254 -6786 497834 30338
rect 504814 704838 505394 705770
rect 504814 704602 504986 704838
rect 505222 704602 505394 704838
rect 504814 704518 505394 704602
rect 504814 704282 504986 704518
rect 505222 704282 505394 704518
rect 504814 686454 505394 704282
rect 504814 686218 504986 686454
rect 505222 686218 505394 686454
rect 504814 686134 505394 686218
rect 504814 685898 504986 686134
rect 505222 685898 505394 686134
rect 504814 650454 505394 685898
rect 504814 650218 504986 650454
rect 505222 650218 505394 650454
rect 504814 650134 505394 650218
rect 504814 649898 504986 650134
rect 505222 649898 505394 650134
rect 504814 614454 505394 649898
rect 504814 614218 504986 614454
rect 505222 614218 505394 614454
rect 504814 614134 505394 614218
rect 504814 613898 504986 614134
rect 505222 613898 505394 614134
rect 504814 578454 505394 613898
rect 504814 578218 504986 578454
rect 505222 578218 505394 578454
rect 504814 578134 505394 578218
rect 504814 577898 504986 578134
rect 505222 577898 505394 578134
rect 504814 542454 505394 577898
rect 504814 542218 504986 542454
rect 505222 542218 505394 542454
rect 504814 542134 505394 542218
rect 504814 541898 504986 542134
rect 505222 541898 505394 542134
rect 504814 506454 505394 541898
rect 504814 506218 504986 506454
rect 505222 506218 505394 506454
rect 504814 506134 505394 506218
rect 504814 505898 504986 506134
rect 505222 505898 505394 506134
rect 504814 470454 505394 505898
rect 504814 470218 504986 470454
rect 505222 470218 505394 470454
rect 504814 470134 505394 470218
rect 504814 469898 504986 470134
rect 505222 469898 505394 470134
rect 504814 434454 505394 469898
rect 504814 434218 504986 434454
rect 505222 434218 505394 434454
rect 504814 434134 505394 434218
rect 504814 433898 504986 434134
rect 505222 433898 505394 434134
rect 504814 398454 505394 433898
rect 504814 398218 504986 398454
rect 505222 398218 505394 398454
rect 504814 398134 505394 398218
rect 504814 397898 504986 398134
rect 505222 397898 505394 398134
rect 504814 362454 505394 397898
rect 504814 362218 504986 362454
rect 505222 362218 505394 362454
rect 504814 362134 505394 362218
rect 504814 361898 504986 362134
rect 505222 361898 505394 362134
rect 504814 326454 505394 361898
rect 504814 326218 504986 326454
rect 505222 326218 505394 326454
rect 504814 326134 505394 326218
rect 504814 325898 504986 326134
rect 505222 325898 505394 326134
rect 504814 290454 505394 325898
rect 504814 290218 504986 290454
rect 505222 290218 505394 290454
rect 504814 290134 505394 290218
rect 504814 289898 504986 290134
rect 505222 289898 505394 290134
rect 504814 254454 505394 289898
rect 504814 254218 504986 254454
rect 505222 254218 505394 254454
rect 504814 254134 505394 254218
rect 504814 253898 504986 254134
rect 505222 253898 505394 254134
rect 504814 218454 505394 253898
rect 504814 218218 504986 218454
rect 505222 218218 505394 218454
rect 504814 218134 505394 218218
rect 504814 217898 504986 218134
rect 505222 217898 505394 218134
rect 504814 182454 505394 217898
rect 504814 182218 504986 182454
rect 505222 182218 505394 182454
rect 504814 182134 505394 182218
rect 504814 181898 504986 182134
rect 505222 181898 505394 182134
rect 504814 146454 505394 181898
rect 504814 146218 504986 146454
rect 505222 146218 505394 146454
rect 504814 146134 505394 146218
rect 504814 145898 504986 146134
rect 505222 145898 505394 146134
rect 504814 110454 505394 145898
rect 504814 110218 504986 110454
rect 505222 110218 505394 110454
rect 504814 110134 505394 110218
rect 504814 109898 504986 110134
rect 505222 109898 505394 110134
rect 504814 74454 505394 109898
rect 504814 74218 504986 74454
rect 505222 74218 505394 74454
rect 504814 74134 505394 74218
rect 504814 73898 504986 74134
rect 505222 73898 505394 74134
rect 504814 38454 505394 73898
rect 504814 38218 504986 38454
rect 505222 38218 505394 38454
rect 504814 38134 505394 38218
rect 504814 37898 504986 38134
rect 505222 37898 505394 38134
rect 504814 2454 505394 37898
rect 504814 2218 504986 2454
rect 505222 2218 505394 2454
rect 504814 2134 505394 2218
rect 504814 1898 504986 2134
rect 505222 1898 505394 2134
rect 504814 -346 505394 1898
rect 504814 -582 504986 -346
rect 505222 -582 505394 -346
rect 504814 -666 505394 -582
rect 504814 -902 504986 -666
rect 505222 -902 505394 -666
rect 504814 -1834 505394 -902
rect 508294 689934 508874 706122
rect 508294 689698 508466 689934
rect 508702 689698 508874 689934
rect 508294 689614 508874 689698
rect 508294 689378 508466 689614
rect 508702 689378 508874 689614
rect 508294 653934 508874 689378
rect 508294 653698 508466 653934
rect 508702 653698 508874 653934
rect 508294 653614 508874 653698
rect 508294 653378 508466 653614
rect 508702 653378 508874 653614
rect 508294 617934 508874 653378
rect 508294 617698 508466 617934
rect 508702 617698 508874 617934
rect 508294 617614 508874 617698
rect 508294 617378 508466 617614
rect 508702 617378 508874 617614
rect 508294 581934 508874 617378
rect 508294 581698 508466 581934
rect 508702 581698 508874 581934
rect 508294 581614 508874 581698
rect 508294 581378 508466 581614
rect 508702 581378 508874 581614
rect 508294 545934 508874 581378
rect 508294 545698 508466 545934
rect 508702 545698 508874 545934
rect 508294 545614 508874 545698
rect 508294 545378 508466 545614
rect 508702 545378 508874 545614
rect 508294 509934 508874 545378
rect 508294 509698 508466 509934
rect 508702 509698 508874 509934
rect 508294 509614 508874 509698
rect 508294 509378 508466 509614
rect 508702 509378 508874 509614
rect 508294 473934 508874 509378
rect 508294 473698 508466 473934
rect 508702 473698 508874 473934
rect 508294 473614 508874 473698
rect 508294 473378 508466 473614
rect 508702 473378 508874 473614
rect 508294 437934 508874 473378
rect 508294 437698 508466 437934
rect 508702 437698 508874 437934
rect 508294 437614 508874 437698
rect 508294 437378 508466 437614
rect 508702 437378 508874 437614
rect 508294 401934 508874 437378
rect 508294 401698 508466 401934
rect 508702 401698 508874 401934
rect 508294 401614 508874 401698
rect 508294 401378 508466 401614
rect 508702 401378 508874 401614
rect 508294 365934 508874 401378
rect 508294 365698 508466 365934
rect 508702 365698 508874 365934
rect 508294 365614 508874 365698
rect 508294 365378 508466 365614
rect 508702 365378 508874 365614
rect 508294 329934 508874 365378
rect 508294 329698 508466 329934
rect 508702 329698 508874 329934
rect 508294 329614 508874 329698
rect 508294 329378 508466 329614
rect 508702 329378 508874 329614
rect 508294 293934 508874 329378
rect 508294 293698 508466 293934
rect 508702 293698 508874 293934
rect 508294 293614 508874 293698
rect 508294 293378 508466 293614
rect 508702 293378 508874 293614
rect 508294 257934 508874 293378
rect 508294 257698 508466 257934
rect 508702 257698 508874 257934
rect 508294 257614 508874 257698
rect 508294 257378 508466 257614
rect 508702 257378 508874 257614
rect 508294 221934 508874 257378
rect 508294 221698 508466 221934
rect 508702 221698 508874 221934
rect 508294 221614 508874 221698
rect 508294 221378 508466 221614
rect 508702 221378 508874 221614
rect 508294 185934 508874 221378
rect 508294 185698 508466 185934
rect 508702 185698 508874 185934
rect 508294 185614 508874 185698
rect 508294 185378 508466 185614
rect 508702 185378 508874 185614
rect 508294 149934 508874 185378
rect 508294 149698 508466 149934
rect 508702 149698 508874 149934
rect 508294 149614 508874 149698
rect 508294 149378 508466 149614
rect 508702 149378 508874 149614
rect 508294 113934 508874 149378
rect 508294 113698 508466 113934
rect 508702 113698 508874 113934
rect 508294 113614 508874 113698
rect 508294 113378 508466 113614
rect 508702 113378 508874 113614
rect 508294 77934 508874 113378
rect 508294 77698 508466 77934
rect 508702 77698 508874 77934
rect 508294 77614 508874 77698
rect 508294 77378 508466 77614
rect 508702 77378 508874 77614
rect 508294 41934 508874 77378
rect 508294 41698 508466 41934
rect 508702 41698 508874 41934
rect 508294 41614 508874 41698
rect 508294 41378 508466 41614
rect 508702 41378 508874 41614
rect 508294 5934 508874 41378
rect 508294 5698 508466 5934
rect 508702 5698 508874 5934
rect 508294 5614 508874 5698
rect 508294 5378 508466 5614
rect 508702 5378 508874 5614
rect 508294 -2186 508874 5378
rect 508294 -2422 508466 -2186
rect 508702 -2422 508874 -2186
rect 508294 -2506 508874 -2422
rect 508294 -2742 508466 -2506
rect 508702 -2742 508874 -2506
rect 508294 -3674 508874 -2742
rect 511774 693414 512354 707962
rect 511774 693178 511946 693414
rect 512182 693178 512354 693414
rect 511774 693094 512354 693178
rect 511774 692858 511946 693094
rect 512182 692858 512354 693094
rect 511774 657414 512354 692858
rect 511774 657178 511946 657414
rect 512182 657178 512354 657414
rect 511774 657094 512354 657178
rect 511774 656858 511946 657094
rect 512182 656858 512354 657094
rect 511774 621414 512354 656858
rect 511774 621178 511946 621414
rect 512182 621178 512354 621414
rect 511774 621094 512354 621178
rect 511774 620858 511946 621094
rect 512182 620858 512354 621094
rect 511774 585414 512354 620858
rect 511774 585178 511946 585414
rect 512182 585178 512354 585414
rect 511774 585094 512354 585178
rect 511774 584858 511946 585094
rect 512182 584858 512354 585094
rect 511774 549414 512354 584858
rect 511774 549178 511946 549414
rect 512182 549178 512354 549414
rect 511774 549094 512354 549178
rect 511774 548858 511946 549094
rect 512182 548858 512354 549094
rect 511774 513414 512354 548858
rect 511774 513178 511946 513414
rect 512182 513178 512354 513414
rect 511774 513094 512354 513178
rect 511774 512858 511946 513094
rect 512182 512858 512354 513094
rect 511774 477414 512354 512858
rect 511774 477178 511946 477414
rect 512182 477178 512354 477414
rect 511774 477094 512354 477178
rect 511774 476858 511946 477094
rect 512182 476858 512354 477094
rect 511774 441414 512354 476858
rect 511774 441178 511946 441414
rect 512182 441178 512354 441414
rect 511774 441094 512354 441178
rect 511774 440858 511946 441094
rect 512182 440858 512354 441094
rect 511774 405414 512354 440858
rect 511774 405178 511946 405414
rect 512182 405178 512354 405414
rect 511774 405094 512354 405178
rect 511774 404858 511946 405094
rect 512182 404858 512354 405094
rect 511774 369414 512354 404858
rect 511774 369178 511946 369414
rect 512182 369178 512354 369414
rect 511774 369094 512354 369178
rect 511774 368858 511946 369094
rect 512182 368858 512354 369094
rect 511774 333414 512354 368858
rect 511774 333178 511946 333414
rect 512182 333178 512354 333414
rect 511774 333094 512354 333178
rect 511774 332858 511946 333094
rect 512182 332858 512354 333094
rect 511774 297414 512354 332858
rect 511774 297178 511946 297414
rect 512182 297178 512354 297414
rect 511774 297094 512354 297178
rect 511774 296858 511946 297094
rect 512182 296858 512354 297094
rect 511774 261414 512354 296858
rect 511774 261178 511946 261414
rect 512182 261178 512354 261414
rect 511774 261094 512354 261178
rect 511774 260858 511946 261094
rect 512182 260858 512354 261094
rect 511774 225414 512354 260858
rect 511774 225178 511946 225414
rect 512182 225178 512354 225414
rect 511774 225094 512354 225178
rect 511774 224858 511946 225094
rect 512182 224858 512354 225094
rect 511774 189414 512354 224858
rect 511774 189178 511946 189414
rect 512182 189178 512354 189414
rect 511774 189094 512354 189178
rect 511774 188858 511946 189094
rect 512182 188858 512354 189094
rect 511774 153414 512354 188858
rect 511774 153178 511946 153414
rect 512182 153178 512354 153414
rect 511774 153094 512354 153178
rect 511774 152858 511946 153094
rect 512182 152858 512354 153094
rect 511774 117414 512354 152858
rect 511774 117178 511946 117414
rect 512182 117178 512354 117414
rect 511774 117094 512354 117178
rect 511774 116858 511946 117094
rect 512182 116858 512354 117094
rect 511774 81414 512354 116858
rect 511774 81178 511946 81414
rect 512182 81178 512354 81414
rect 511774 81094 512354 81178
rect 511774 80858 511946 81094
rect 512182 80858 512354 81094
rect 511774 45414 512354 80858
rect 511774 45178 511946 45414
rect 512182 45178 512354 45414
rect 511774 45094 512354 45178
rect 511774 44858 511946 45094
rect 512182 44858 512354 45094
rect 511774 9414 512354 44858
rect 511774 9178 511946 9414
rect 512182 9178 512354 9414
rect 511774 9094 512354 9178
rect 511774 8858 511946 9094
rect 512182 8858 512354 9094
rect 511774 -4026 512354 8858
rect 511774 -4262 511946 -4026
rect 512182 -4262 512354 -4026
rect 511774 -4346 512354 -4262
rect 511774 -4582 511946 -4346
rect 512182 -4582 512354 -4346
rect 511774 -5514 512354 -4582
rect 515254 696894 515834 709802
rect 533254 711278 533834 711290
rect 533254 711042 533426 711278
rect 533662 711042 533834 711278
rect 533254 710958 533834 711042
rect 533254 710722 533426 710958
rect 533662 710722 533834 710958
rect 529774 709438 530354 709450
rect 529774 709202 529946 709438
rect 530182 709202 530354 709438
rect 529774 709118 530354 709202
rect 529774 708882 529946 709118
rect 530182 708882 530354 709118
rect 526294 707598 526874 707610
rect 526294 707362 526466 707598
rect 526702 707362 526874 707598
rect 526294 707278 526874 707362
rect 526294 707042 526466 707278
rect 526702 707042 526874 707278
rect 515254 696658 515426 696894
rect 515662 696658 515834 696894
rect 515254 696574 515834 696658
rect 515254 696338 515426 696574
rect 515662 696338 515834 696574
rect 515254 660894 515834 696338
rect 515254 660658 515426 660894
rect 515662 660658 515834 660894
rect 515254 660574 515834 660658
rect 515254 660338 515426 660574
rect 515662 660338 515834 660574
rect 515254 624894 515834 660338
rect 515254 624658 515426 624894
rect 515662 624658 515834 624894
rect 515254 624574 515834 624658
rect 515254 624338 515426 624574
rect 515662 624338 515834 624574
rect 515254 588894 515834 624338
rect 515254 588658 515426 588894
rect 515662 588658 515834 588894
rect 515254 588574 515834 588658
rect 515254 588338 515426 588574
rect 515662 588338 515834 588574
rect 515254 552894 515834 588338
rect 515254 552658 515426 552894
rect 515662 552658 515834 552894
rect 515254 552574 515834 552658
rect 515254 552338 515426 552574
rect 515662 552338 515834 552574
rect 515254 516894 515834 552338
rect 515254 516658 515426 516894
rect 515662 516658 515834 516894
rect 515254 516574 515834 516658
rect 515254 516338 515426 516574
rect 515662 516338 515834 516574
rect 515254 480894 515834 516338
rect 515254 480658 515426 480894
rect 515662 480658 515834 480894
rect 515254 480574 515834 480658
rect 515254 480338 515426 480574
rect 515662 480338 515834 480574
rect 515254 444894 515834 480338
rect 515254 444658 515426 444894
rect 515662 444658 515834 444894
rect 515254 444574 515834 444658
rect 515254 444338 515426 444574
rect 515662 444338 515834 444574
rect 515254 408894 515834 444338
rect 515254 408658 515426 408894
rect 515662 408658 515834 408894
rect 515254 408574 515834 408658
rect 515254 408338 515426 408574
rect 515662 408338 515834 408574
rect 515254 372894 515834 408338
rect 515254 372658 515426 372894
rect 515662 372658 515834 372894
rect 515254 372574 515834 372658
rect 515254 372338 515426 372574
rect 515662 372338 515834 372574
rect 515254 336894 515834 372338
rect 515254 336658 515426 336894
rect 515662 336658 515834 336894
rect 515254 336574 515834 336658
rect 515254 336338 515426 336574
rect 515662 336338 515834 336574
rect 515254 300894 515834 336338
rect 515254 300658 515426 300894
rect 515662 300658 515834 300894
rect 515254 300574 515834 300658
rect 515254 300338 515426 300574
rect 515662 300338 515834 300574
rect 515254 264894 515834 300338
rect 515254 264658 515426 264894
rect 515662 264658 515834 264894
rect 515254 264574 515834 264658
rect 515254 264338 515426 264574
rect 515662 264338 515834 264574
rect 515254 228894 515834 264338
rect 515254 228658 515426 228894
rect 515662 228658 515834 228894
rect 515254 228574 515834 228658
rect 515254 228338 515426 228574
rect 515662 228338 515834 228574
rect 515254 192894 515834 228338
rect 515254 192658 515426 192894
rect 515662 192658 515834 192894
rect 515254 192574 515834 192658
rect 515254 192338 515426 192574
rect 515662 192338 515834 192574
rect 515254 156894 515834 192338
rect 515254 156658 515426 156894
rect 515662 156658 515834 156894
rect 515254 156574 515834 156658
rect 515254 156338 515426 156574
rect 515662 156338 515834 156574
rect 515254 120894 515834 156338
rect 515254 120658 515426 120894
rect 515662 120658 515834 120894
rect 515254 120574 515834 120658
rect 515254 120338 515426 120574
rect 515662 120338 515834 120574
rect 515254 84894 515834 120338
rect 515254 84658 515426 84894
rect 515662 84658 515834 84894
rect 515254 84574 515834 84658
rect 515254 84338 515426 84574
rect 515662 84338 515834 84574
rect 515254 48894 515834 84338
rect 515254 48658 515426 48894
rect 515662 48658 515834 48894
rect 515254 48574 515834 48658
rect 515254 48338 515426 48574
rect 515662 48338 515834 48574
rect 515254 12894 515834 48338
rect 515254 12658 515426 12894
rect 515662 12658 515834 12894
rect 515254 12574 515834 12658
rect 515254 12338 515426 12574
rect 515662 12338 515834 12574
rect 497254 -7022 497426 -6786
rect 497662 -7022 497834 -6786
rect 497254 -7106 497834 -7022
rect 497254 -7342 497426 -7106
rect 497662 -7342 497834 -7106
rect 497254 -7354 497834 -7342
rect 515254 -5866 515834 12338
rect 522814 705758 523394 705770
rect 522814 705522 522986 705758
rect 523222 705522 523394 705758
rect 522814 705438 523394 705522
rect 522814 705202 522986 705438
rect 523222 705202 523394 705438
rect 522814 668454 523394 705202
rect 522814 668218 522986 668454
rect 523222 668218 523394 668454
rect 522814 668134 523394 668218
rect 522814 667898 522986 668134
rect 523222 667898 523394 668134
rect 522814 632454 523394 667898
rect 522814 632218 522986 632454
rect 523222 632218 523394 632454
rect 522814 632134 523394 632218
rect 522814 631898 522986 632134
rect 523222 631898 523394 632134
rect 522814 596454 523394 631898
rect 522814 596218 522986 596454
rect 523222 596218 523394 596454
rect 522814 596134 523394 596218
rect 522814 595898 522986 596134
rect 523222 595898 523394 596134
rect 522814 560454 523394 595898
rect 522814 560218 522986 560454
rect 523222 560218 523394 560454
rect 522814 560134 523394 560218
rect 522814 559898 522986 560134
rect 523222 559898 523394 560134
rect 522814 524454 523394 559898
rect 522814 524218 522986 524454
rect 523222 524218 523394 524454
rect 522814 524134 523394 524218
rect 522814 523898 522986 524134
rect 523222 523898 523394 524134
rect 522814 488454 523394 523898
rect 522814 488218 522986 488454
rect 523222 488218 523394 488454
rect 522814 488134 523394 488218
rect 522814 487898 522986 488134
rect 523222 487898 523394 488134
rect 522814 452454 523394 487898
rect 522814 452218 522986 452454
rect 523222 452218 523394 452454
rect 522814 452134 523394 452218
rect 522814 451898 522986 452134
rect 523222 451898 523394 452134
rect 522814 416454 523394 451898
rect 522814 416218 522986 416454
rect 523222 416218 523394 416454
rect 522814 416134 523394 416218
rect 522814 415898 522986 416134
rect 523222 415898 523394 416134
rect 522814 380454 523394 415898
rect 522814 380218 522986 380454
rect 523222 380218 523394 380454
rect 522814 380134 523394 380218
rect 522814 379898 522986 380134
rect 523222 379898 523394 380134
rect 522814 344454 523394 379898
rect 522814 344218 522986 344454
rect 523222 344218 523394 344454
rect 522814 344134 523394 344218
rect 522814 343898 522986 344134
rect 523222 343898 523394 344134
rect 522814 308454 523394 343898
rect 522814 308218 522986 308454
rect 523222 308218 523394 308454
rect 522814 308134 523394 308218
rect 522814 307898 522986 308134
rect 523222 307898 523394 308134
rect 522814 272454 523394 307898
rect 522814 272218 522986 272454
rect 523222 272218 523394 272454
rect 522814 272134 523394 272218
rect 522814 271898 522986 272134
rect 523222 271898 523394 272134
rect 522814 236454 523394 271898
rect 522814 236218 522986 236454
rect 523222 236218 523394 236454
rect 522814 236134 523394 236218
rect 522814 235898 522986 236134
rect 523222 235898 523394 236134
rect 522814 200454 523394 235898
rect 522814 200218 522986 200454
rect 523222 200218 523394 200454
rect 522814 200134 523394 200218
rect 522814 199898 522986 200134
rect 523222 199898 523394 200134
rect 522814 164454 523394 199898
rect 522814 164218 522986 164454
rect 523222 164218 523394 164454
rect 522814 164134 523394 164218
rect 522814 163898 522986 164134
rect 523222 163898 523394 164134
rect 522814 128454 523394 163898
rect 522814 128218 522986 128454
rect 523222 128218 523394 128454
rect 522814 128134 523394 128218
rect 522814 127898 522986 128134
rect 523222 127898 523394 128134
rect 522814 92454 523394 127898
rect 522814 92218 522986 92454
rect 523222 92218 523394 92454
rect 522814 92134 523394 92218
rect 522814 91898 522986 92134
rect 523222 91898 523394 92134
rect 522814 56454 523394 91898
rect 522814 56218 522986 56454
rect 523222 56218 523394 56454
rect 522814 56134 523394 56218
rect 522814 55898 522986 56134
rect 523222 55898 523394 56134
rect 522814 20454 523394 55898
rect 522814 20218 522986 20454
rect 523222 20218 523394 20454
rect 522814 20134 523394 20218
rect 522814 19898 522986 20134
rect 523222 19898 523394 20134
rect 522814 -1266 523394 19898
rect 522814 -1502 522986 -1266
rect 523222 -1502 523394 -1266
rect 522814 -1586 523394 -1502
rect 522814 -1822 522986 -1586
rect 523222 -1822 523394 -1586
rect 522814 -1834 523394 -1822
rect 526294 671934 526874 707042
rect 526294 671698 526466 671934
rect 526702 671698 526874 671934
rect 526294 671614 526874 671698
rect 526294 671378 526466 671614
rect 526702 671378 526874 671614
rect 526294 635934 526874 671378
rect 526294 635698 526466 635934
rect 526702 635698 526874 635934
rect 526294 635614 526874 635698
rect 526294 635378 526466 635614
rect 526702 635378 526874 635614
rect 526294 599934 526874 635378
rect 526294 599698 526466 599934
rect 526702 599698 526874 599934
rect 526294 599614 526874 599698
rect 526294 599378 526466 599614
rect 526702 599378 526874 599614
rect 526294 563934 526874 599378
rect 526294 563698 526466 563934
rect 526702 563698 526874 563934
rect 526294 563614 526874 563698
rect 526294 563378 526466 563614
rect 526702 563378 526874 563614
rect 526294 527934 526874 563378
rect 526294 527698 526466 527934
rect 526702 527698 526874 527934
rect 526294 527614 526874 527698
rect 526294 527378 526466 527614
rect 526702 527378 526874 527614
rect 526294 491934 526874 527378
rect 526294 491698 526466 491934
rect 526702 491698 526874 491934
rect 526294 491614 526874 491698
rect 526294 491378 526466 491614
rect 526702 491378 526874 491614
rect 526294 455934 526874 491378
rect 526294 455698 526466 455934
rect 526702 455698 526874 455934
rect 526294 455614 526874 455698
rect 526294 455378 526466 455614
rect 526702 455378 526874 455614
rect 526294 419934 526874 455378
rect 526294 419698 526466 419934
rect 526702 419698 526874 419934
rect 526294 419614 526874 419698
rect 526294 419378 526466 419614
rect 526702 419378 526874 419614
rect 526294 383934 526874 419378
rect 526294 383698 526466 383934
rect 526702 383698 526874 383934
rect 526294 383614 526874 383698
rect 526294 383378 526466 383614
rect 526702 383378 526874 383614
rect 526294 347934 526874 383378
rect 526294 347698 526466 347934
rect 526702 347698 526874 347934
rect 526294 347614 526874 347698
rect 526294 347378 526466 347614
rect 526702 347378 526874 347614
rect 526294 311934 526874 347378
rect 526294 311698 526466 311934
rect 526702 311698 526874 311934
rect 526294 311614 526874 311698
rect 526294 311378 526466 311614
rect 526702 311378 526874 311614
rect 526294 275934 526874 311378
rect 526294 275698 526466 275934
rect 526702 275698 526874 275934
rect 526294 275614 526874 275698
rect 526294 275378 526466 275614
rect 526702 275378 526874 275614
rect 526294 239934 526874 275378
rect 526294 239698 526466 239934
rect 526702 239698 526874 239934
rect 526294 239614 526874 239698
rect 526294 239378 526466 239614
rect 526702 239378 526874 239614
rect 526294 203934 526874 239378
rect 526294 203698 526466 203934
rect 526702 203698 526874 203934
rect 526294 203614 526874 203698
rect 526294 203378 526466 203614
rect 526702 203378 526874 203614
rect 526294 167934 526874 203378
rect 526294 167698 526466 167934
rect 526702 167698 526874 167934
rect 526294 167614 526874 167698
rect 526294 167378 526466 167614
rect 526702 167378 526874 167614
rect 526294 131934 526874 167378
rect 526294 131698 526466 131934
rect 526702 131698 526874 131934
rect 526294 131614 526874 131698
rect 526294 131378 526466 131614
rect 526702 131378 526874 131614
rect 526294 95934 526874 131378
rect 526294 95698 526466 95934
rect 526702 95698 526874 95934
rect 526294 95614 526874 95698
rect 526294 95378 526466 95614
rect 526702 95378 526874 95614
rect 526294 59934 526874 95378
rect 526294 59698 526466 59934
rect 526702 59698 526874 59934
rect 526294 59614 526874 59698
rect 526294 59378 526466 59614
rect 526702 59378 526874 59614
rect 526294 23934 526874 59378
rect 526294 23698 526466 23934
rect 526702 23698 526874 23934
rect 526294 23614 526874 23698
rect 526294 23378 526466 23614
rect 526702 23378 526874 23614
rect 526294 -3106 526874 23378
rect 526294 -3342 526466 -3106
rect 526702 -3342 526874 -3106
rect 526294 -3426 526874 -3342
rect 526294 -3662 526466 -3426
rect 526702 -3662 526874 -3426
rect 526294 -3674 526874 -3662
rect 529774 675414 530354 708882
rect 529774 675178 529946 675414
rect 530182 675178 530354 675414
rect 529774 675094 530354 675178
rect 529774 674858 529946 675094
rect 530182 674858 530354 675094
rect 529774 639414 530354 674858
rect 529774 639178 529946 639414
rect 530182 639178 530354 639414
rect 529774 639094 530354 639178
rect 529774 638858 529946 639094
rect 530182 638858 530354 639094
rect 529774 603414 530354 638858
rect 529774 603178 529946 603414
rect 530182 603178 530354 603414
rect 529774 603094 530354 603178
rect 529774 602858 529946 603094
rect 530182 602858 530354 603094
rect 529774 567414 530354 602858
rect 529774 567178 529946 567414
rect 530182 567178 530354 567414
rect 529774 567094 530354 567178
rect 529774 566858 529946 567094
rect 530182 566858 530354 567094
rect 529774 531414 530354 566858
rect 529774 531178 529946 531414
rect 530182 531178 530354 531414
rect 529774 531094 530354 531178
rect 529774 530858 529946 531094
rect 530182 530858 530354 531094
rect 529774 495414 530354 530858
rect 529774 495178 529946 495414
rect 530182 495178 530354 495414
rect 529774 495094 530354 495178
rect 529774 494858 529946 495094
rect 530182 494858 530354 495094
rect 529774 459414 530354 494858
rect 529774 459178 529946 459414
rect 530182 459178 530354 459414
rect 529774 459094 530354 459178
rect 529774 458858 529946 459094
rect 530182 458858 530354 459094
rect 529774 423414 530354 458858
rect 529774 423178 529946 423414
rect 530182 423178 530354 423414
rect 529774 423094 530354 423178
rect 529774 422858 529946 423094
rect 530182 422858 530354 423094
rect 529774 387414 530354 422858
rect 529774 387178 529946 387414
rect 530182 387178 530354 387414
rect 529774 387094 530354 387178
rect 529774 386858 529946 387094
rect 530182 386858 530354 387094
rect 529774 351414 530354 386858
rect 529774 351178 529946 351414
rect 530182 351178 530354 351414
rect 529774 351094 530354 351178
rect 529774 350858 529946 351094
rect 530182 350858 530354 351094
rect 529774 315414 530354 350858
rect 529774 315178 529946 315414
rect 530182 315178 530354 315414
rect 529774 315094 530354 315178
rect 529774 314858 529946 315094
rect 530182 314858 530354 315094
rect 529774 279414 530354 314858
rect 529774 279178 529946 279414
rect 530182 279178 530354 279414
rect 529774 279094 530354 279178
rect 529774 278858 529946 279094
rect 530182 278858 530354 279094
rect 529774 243414 530354 278858
rect 529774 243178 529946 243414
rect 530182 243178 530354 243414
rect 529774 243094 530354 243178
rect 529774 242858 529946 243094
rect 530182 242858 530354 243094
rect 529774 207414 530354 242858
rect 529774 207178 529946 207414
rect 530182 207178 530354 207414
rect 529774 207094 530354 207178
rect 529774 206858 529946 207094
rect 530182 206858 530354 207094
rect 529774 171414 530354 206858
rect 529774 171178 529946 171414
rect 530182 171178 530354 171414
rect 529774 171094 530354 171178
rect 529774 170858 529946 171094
rect 530182 170858 530354 171094
rect 529774 135414 530354 170858
rect 529774 135178 529946 135414
rect 530182 135178 530354 135414
rect 529774 135094 530354 135178
rect 529774 134858 529946 135094
rect 530182 134858 530354 135094
rect 529774 99414 530354 134858
rect 529774 99178 529946 99414
rect 530182 99178 530354 99414
rect 529774 99094 530354 99178
rect 529774 98858 529946 99094
rect 530182 98858 530354 99094
rect 529774 63414 530354 98858
rect 529774 63178 529946 63414
rect 530182 63178 530354 63414
rect 529774 63094 530354 63178
rect 529774 62858 529946 63094
rect 530182 62858 530354 63094
rect 529774 27414 530354 62858
rect 529774 27178 529946 27414
rect 530182 27178 530354 27414
rect 529774 27094 530354 27178
rect 529774 26858 529946 27094
rect 530182 26858 530354 27094
rect 529774 -4946 530354 26858
rect 529774 -5182 529946 -4946
rect 530182 -5182 530354 -4946
rect 529774 -5266 530354 -5182
rect 529774 -5502 529946 -5266
rect 530182 -5502 530354 -5266
rect 529774 -5514 530354 -5502
rect 533254 678894 533834 710722
rect 551254 710358 551834 711290
rect 551254 710122 551426 710358
rect 551662 710122 551834 710358
rect 551254 710038 551834 710122
rect 551254 709802 551426 710038
rect 551662 709802 551834 710038
rect 547774 708518 548354 709450
rect 547774 708282 547946 708518
rect 548182 708282 548354 708518
rect 547774 708198 548354 708282
rect 547774 707962 547946 708198
rect 548182 707962 548354 708198
rect 544294 706678 544874 707610
rect 544294 706442 544466 706678
rect 544702 706442 544874 706678
rect 544294 706358 544874 706442
rect 544294 706122 544466 706358
rect 544702 706122 544874 706358
rect 533254 678658 533426 678894
rect 533662 678658 533834 678894
rect 533254 678574 533834 678658
rect 533254 678338 533426 678574
rect 533662 678338 533834 678574
rect 533254 642894 533834 678338
rect 533254 642658 533426 642894
rect 533662 642658 533834 642894
rect 533254 642574 533834 642658
rect 533254 642338 533426 642574
rect 533662 642338 533834 642574
rect 533254 606894 533834 642338
rect 533254 606658 533426 606894
rect 533662 606658 533834 606894
rect 533254 606574 533834 606658
rect 533254 606338 533426 606574
rect 533662 606338 533834 606574
rect 533254 570894 533834 606338
rect 533254 570658 533426 570894
rect 533662 570658 533834 570894
rect 533254 570574 533834 570658
rect 533254 570338 533426 570574
rect 533662 570338 533834 570574
rect 533254 534894 533834 570338
rect 533254 534658 533426 534894
rect 533662 534658 533834 534894
rect 533254 534574 533834 534658
rect 533254 534338 533426 534574
rect 533662 534338 533834 534574
rect 533254 498894 533834 534338
rect 533254 498658 533426 498894
rect 533662 498658 533834 498894
rect 533254 498574 533834 498658
rect 533254 498338 533426 498574
rect 533662 498338 533834 498574
rect 533254 462894 533834 498338
rect 533254 462658 533426 462894
rect 533662 462658 533834 462894
rect 533254 462574 533834 462658
rect 533254 462338 533426 462574
rect 533662 462338 533834 462574
rect 533254 426894 533834 462338
rect 533254 426658 533426 426894
rect 533662 426658 533834 426894
rect 533254 426574 533834 426658
rect 533254 426338 533426 426574
rect 533662 426338 533834 426574
rect 533254 390894 533834 426338
rect 533254 390658 533426 390894
rect 533662 390658 533834 390894
rect 533254 390574 533834 390658
rect 533254 390338 533426 390574
rect 533662 390338 533834 390574
rect 533254 354894 533834 390338
rect 533254 354658 533426 354894
rect 533662 354658 533834 354894
rect 533254 354574 533834 354658
rect 533254 354338 533426 354574
rect 533662 354338 533834 354574
rect 533254 318894 533834 354338
rect 533254 318658 533426 318894
rect 533662 318658 533834 318894
rect 533254 318574 533834 318658
rect 533254 318338 533426 318574
rect 533662 318338 533834 318574
rect 533254 282894 533834 318338
rect 533254 282658 533426 282894
rect 533662 282658 533834 282894
rect 533254 282574 533834 282658
rect 533254 282338 533426 282574
rect 533662 282338 533834 282574
rect 533254 246894 533834 282338
rect 533254 246658 533426 246894
rect 533662 246658 533834 246894
rect 533254 246574 533834 246658
rect 533254 246338 533426 246574
rect 533662 246338 533834 246574
rect 533254 210894 533834 246338
rect 533254 210658 533426 210894
rect 533662 210658 533834 210894
rect 533254 210574 533834 210658
rect 533254 210338 533426 210574
rect 533662 210338 533834 210574
rect 533254 174894 533834 210338
rect 533254 174658 533426 174894
rect 533662 174658 533834 174894
rect 533254 174574 533834 174658
rect 533254 174338 533426 174574
rect 533662 174338 533834 174574
rect 533254 138894 533834 174338
rect 533254 138658 533426 138894
rect 533662 138658 533834 138894
rect 533254 138574 533834 138658
rect 533254 138338 533426 138574
rect 533662 138338 533834 138574
rect 533254 102894 533834 138338
rect 533254 102658 533426 102894
rect 533662 102658 533834 102894
rect 533254 102574 533834 102658
rect 533254 102338 533426 102574
rect 533662 102338 533834 102574
rect 533254 66894 533834 102338
rect 533254 66658 533426 66894
rect 533662 66658 533834 66894
rect 533254 66574 533834 66658
rect 533254 66338 533426 66574
rect 533662 66338 533834 66574
rect 533254 30894 533834 66338
rect 533254 30658 533426 30894
rect 533662 30658 533834 30894
rect 533254 30574 533834 30658
rect 533254 30338 533426 30574
rect 533662 30338 533834 30574
rect 515254 -6102 515426 -5866
rect 515662 -6102 515834 -5866
rect 515254 -6186 515834 -6102
rect 515254 -6422 515426 -6186
rect 515662 -6422 515834 -6186
rect 515254 -7354 515834 -6422
rect 533254 -6786 533834 30338
rect 540814 704838 541394 705770
rect 540814 704602 540986 704838
rect 541222 704602 541394 704838
rect 540814 704518 541394 704602
rect 540814 704282 540986 704518
rect 541222 704282 541394 704518
rect 540814 686454 541394 704282
rect 540814 686218 540986 686454
rect 541222 686218 541394 686454
rect 540814 686134 541394 686218
rect 540814 685898 540986 686134
rect 541222 685898 541394 686134
rect 540814 650454 541394 685898
rect 540814 650218 540986 650454
rect 541222 650218 541394 650454
rect 540814 650134 541394 650218
rect 540814 649898 540986 650134
rect 541222 649898 541394 650134
rect 540814 614454 541394 649898
rect 540814 614218 540986 614454
rect 541222 614218 541394 614454
rect 540814 614134 541394 614218
rect 540814 613898 540986 614134
rect 541222 613898 541394 614134
rect 540814 578454 541394 613898
rect 540814 578218 540986 578454
rect 541222 578218 541394 578454
rect 540814 578134 541394 578218
rect 540814 577898 540986 578134
rect 541222 577898 541394 578134
rect 540814 542454 541394 577898
rect 540814 542218 540986 542454
rect 541222 542218 541394 542454
rect 540814 542134 541394 542218
rect 540814 541898 540986 542134
rect 541222 541898 541394 542134
rect 540814 506454 541394 541898
rect 540814 506218 540986 506454
rect 541222 506218 541394 506454
rect 540814 506134 541394 506218
rect 540814 505898 540986 506134
rect 541222 505898 541394 506134
rect 540814 470454 541394 505898
rect 540814 470218 540986 470454
rect 541222 470218 541394 470454
rect 540814 470134 541394 470218
rect 540814 469898 540986 470134
rect 541222 469898 541394 470134
rect 540814 434454 541394 469898
rect 540814 434218 540986 434454
rect 541222 434218 541394 434454
rect 540814 434134 541394 434218
rect 540814 433898 540986 434134
rect 541222 433898 541394 434134
rect 540814 398454 541394 433898
rect 540814 398218 540986 398454
rect 541222 398218 541394 398454
rect 540814 398134 541394 398218
rect 540814 397898 540986 398134
rect 541222 397898 541394 398134
rect 540814 362454 541394 397898
rect 540814 362218 540986 362454
rect 541222 362218 541394 362454
rect 540814 362134 541394 362218
rect 540814 361898 540986 362134
rect 541222 361898 541394 362134
rect 540814 326454 541394 361898
rect 540814 326218 540986 326454
rect 541222 326218 541394 326454
rect 540814 326134 541394 326218
rect 540814 325898 540986 326134
rect 541222 325898 541394 326134
rect 540814 290454 541394 325898
rect 540814 290218 540986 290454
rect 541222 290218 541394 290454
rect 540814 290134 541394 290218
rect 540814 289898 540986 290134
rect 541222 289898 541394 290134
rect 540814 254454 541394 289898
rect 540814 254218 540986 254454
rect 541222 254218 541394 254454
rect 540814 254134 541394 254218
rect 540814 253898 540986 254134
rect 541222 253898 541394 254134
rect 540814 218454 541394 253898
rect 540814 218218 540986 218454
rect 541222 218218 541394 218454
rect 540814 218134 541394 218218
rect 540814 217898 540986 218134
rect 541222 217898 541394 218134
rect 540814 182454 541394 217898
rect 540814 182218 540986 182454
rect 541222 182218 541394 182454
rect 540814 182134 541394 182218
rect 540814 181898 540986 182134
rect 541222 181898 541394 182134
rect 540814 146454 541394 181898
rect 540814 146218 540986 146454
rect 541222 146218 541394 146454
rect 540814 146134 541394 146218
rect 540814 145898 540986 146134
rect 541222 145898 541394 146134
rect 540814 110454 541394 145898
rect 540814 110218 540986 110454
rect 541222 110218 541394 110454
rect 540814 110134 541394 110218
rect 540814 109898 540986 110134
rect 541222 109898 541394 110134
rect 540814 74454 541394 109898
rect 540814 74218 540986 74454
rect 541222 74218 541394 74454
rect 540814 74134 541394 74218
rect 540814 73898 540986 74134
rect 541222 73898 541394 74134
rect 540814 38454 541394 73898
rect 540814 38218 540986 38454
rect 541222 38218 541394 38454
rect 540814 38134 541394 38218
rect 540814 37898 540986 38134
rect 541222 37898 541394 38134
rect 540814 2454 541394 37898
rect 540814 2218 540986 2454
rect 541222 2218 541394 2454
rect 540814 2134 541394 2218
rect 540814 1898 540986 2134
rect 541222 1898 541394 2134
rect 540814 -346 541394 1898
rect 540814 -582 540986 -346
rect 541222 -582 541394 -346
rect 540814 -666 541394 -582
rect 540814 -902 540986 -666
rect 541222 -902 541394 -666
rect 540814 -1834 541394 -902
rect 544294 689934 544874 706122
rect 544294 689698 544466 689934
rect 544702 689698 544874 689934
rect 544294 689614 544874 689698
rect 544294 689378 544466 689614
rect 544702 689378 544874 689614
rect 544294 653934 544874 689378
rect 544294 653698 544466 653934
rect 544702 653698 544874 653934
rect 544294 653614 544874 653698
rect 544294 653378 544466 653614
rect 544702 653378 544874 653614
rect 544294 617934 544874 653378
rect 544294 617698 544466 617934
rect 544702 617698 544874 617934
rect 544294 617614 544874 617698
rect 544294 617378 544466 617614
rect 544702 617378 544874 617614
rect 544294 581934 544874 617378
rect 544294 581698 544466 581934
rect 544702 581698 544874 581934
rect 544294 581614 544874 581698
rect 544294 581378 544466 581614
rect 544702 581378 544874 581614
rect 544294 545934 544874 581378
rect 544294 545698 544466 545934
rect 544702 545698 544874 545934
rect 544294 545614 544874 545698
rect 544294 545378 544466 545614
rect 544702 545378 544874 545614
rect 544294 509934 544874 545378
rect 544294 509698 544466 509934
rect 544702 509698 544874 509934
rect 544294 509614 544874 509698
rect 544294 509378 544466 509614
rect 544702 509378 544874 509614
rect 544294 473934 544874 509378
rect 544294 473698 544466 473934
rect 544702 473698 544874 473934
rect 544294 473614 544874 473698
rect 544294 473378 544466 473614
rect 544702 473378 544874 473614
rect 544294 437934 544874 473378
rect 544294 437698 544466 437934
rect 544702 437698 544874 437934
rect 544294 437614 544874 437698
rect 544294 437378 544466 437614
rect 544702 437378 544874 437614
rect 544294 401934 544874 437378
rect 544294 401698 544466 401934
rect 544702 401698 544874 401934
rect 544294 401614 544874 401698
rect 544294 401378 544466 401614
rect 544702 401378 544874 401614
rect 544294 365934 544874 401378
rect 544294 365698 544466 365934
rect 544702 365698 544874 365934
rect 544294 365614 544874 365698
rect 544294 365378 544466 365614
rect 544702 365378 544874 365614
rect 544294 329934 544874 365378
rect 544294 329698 544466 329934
rect 544702 329698 544874 329934
rect 544294 329614 544874 329698
rect 544294 329378 544466 329614
rect 544702 329378 544874 329614
rect 544294 293934 544874 329378
rect 544294 293698 544466 293934
rect 544702 293698 544874 293934
rect 544294 293614 544874 293698
rect 544294 293378 544466 293614
rect 544702 293378 544874 293614
rect 544294 257934 544874 293378
rect 544294 257698 544466 257934
rect 544702 257698 544874 257934
rect 544294 257614 544874 257698
rect 544294 257378 544466 257614
rect 544702 257378 544874 257614
rect 544294 221934 544874 257378
rect 544294 221698 544466 221934
rect 544702 221698 544874 221934
rect 544294 221614 544874 221698
rect 544294 221378 544466 221614
rect 544702 221378 544874 221614
rect 544294 185934 544874 221378
rect 544294 185698 544466 185934
rect 544702 185698 544874 185934
rect 544294 185614 544874 185698
rect 544294 185378 544466 185614
rect 544702 185378 544874 185614
rect 544294 149934 544874 185378
rect 544294 149698 544466 149934
rect 544702 149698 544874 149934
rect 544294 149614 544874 149698
rect 544294 149378 544466 149614
rect 544702 149378 544874 149614
rect 544294 113934 544874 149378
rect 544294 113698 544466 113934
rect 544702 113698 544874 113934
rect 544294 113614 544874 113698
rect 544294 113378 544466 113614
rect 544702 113378 544874 113614
rect 544294 77934 544874 113378
rect 544294 77698 544466 77934
rect 544702 77698 544874 77934
rect 544294 77614 544874 77698
rect 544294 77378 544466 77614
rect 544702 77378 544874 77614
rect 544294 41934 544874 77378
rect 544294 41698 544466 41934
rect 544702 41698 544874 41934
rect 544294 41614 544874 41698
rect 544294 41378 544466 41614
rect 544702 41378 544874 41614
rect 544294 5934 544874 41378
rect 544294 5698 544466 5934
rect 544702 5698 544874 5934
rect 544294 5614 544874 5698
rect 544294 5378 544466 5614
rect 544702 5378 544874 5614
rect 544294 -2186 544874 5378
rect 544294 -2422 544466 -2186
rect 544702 -2422 544874 -2186
rect 544294 -2506 544874 -2422
rect 544294 -2742 544466 -2506
rect 544702 -2742 544874 -2506
rect 544294 -3674 544874 -2742
rect 547774 693414 548354 707962
rect 547774 693178 547946 693414
rect 548182 693178 548354 693414
rect 547774 693094 548354 693178
rect 547774 692858 547946 693094
rect 548182 692858 548354 693094
rect 547774 657414 548354 692858
rect 547774 657178 547946 657414
rect 548182 657178 548354 657414
rect 547774 657094 548354 657178
rect 547774 656858 547946 657094
rect 548182 656858 548354 657094
rect 547774 621414 548354 656858
rect 547774 621178 547946 621414
rect 548182 621178 548354 621414
rect 547774 621094 548354 621178
rect 547774 620858 547946 621094
rect 548182 620858 548354 621094
rect 547774 585414 548354 620858
rect 547774 585178 547946 585414
rect 548182 585178 548354 585414
rect 547774 585094 548354 585178
rect 547774 584858 547946 585094
rect 548182 584858 548354 585094
rect 547774 549414 548354 584858
rect 547774 549178 547946 549414
rect 548182 549178 548354 549414
rect 547774 549094 548354 549178
rect 547774 548858 547946 549094
rect 548182 548858 548354 549094
rect 547774 513414 548354 548858
rect 547774 513178 547946 513414
rect 548182 513178 548354 513414
rect 547774 513094 548354 513178
rect 547774 512858 547946 513094
rect 548182 512858 548354 513094
rect 547774 477414 548354 512858
rect 547774 477178 547946 477414
rect 548182 477178 548354 477414
rect 547774 477094 548354 477178
rect 547774 476858 547946 477094
rect 548182 476858 548354 477094
rect 547774 441414 548354 476858
rect 547774 441178 547946 441414
rect 548182 441178 548354 441414
rect 547774 441094 548354 441178
rect 547774 440858 547946 441094
rect 548182 440858 548354 441094
rect 547774 405414 548354 440858
rect 547774 405178 547946 405414
rect 548182 405178 548354 405414
rect 547774 405094 548354 405178
rect 547774 404858 547946 405094
rect 548182 404858 548354 405094
rect 547774 369414 548354 404858
rect 547774 369178 547946 369414
rect 548182 369178 548354 369414
rect 547774 369094 548354 369178
rect 547774 368858 547946 369094
rect 548182 368858 548354 369094
rect 547774 333414 548354 368858
rect 547774 333178 547946 333414
rect 548182 333178 548354 333414
rect 547774 333094 548354 333178
rect 547774 332858 547946 333094
rect 548182 332858 548354 333094
rect 547774 297414 548354 332858
rect 547774 297178 547946 297414
rect 548182 297178 548354 297414
rect 547774 297094 548354 297178
rect 547774 296858 547946 297094
rect 548182 296858 548354 297094
rect 547774 261414 548354 296858
rect 547774 261178 547946 261414
rect 548182 261178 548354 261414
rect 547774 261094 548354 261178
rect 547774 260858 547946 261094
rect 548182 260858 548354 261094
rect 547774 225414 548354 260858
rect 547774 225178 547946 225414
rect 548182 225178 548354 225414
rect 547774 225094 548354 225178
rect 547774 224858 547946 225094
rect 548182 224858 548354 225094
rect 547774 189414 548354 224858
rect 547774 189178 547946 189414
rect 548182 189178 548354 189414
rect 547774 189094 548354 189178
rect 547774 188858 547946 189094
rect 548182 188858 548354 189094
rect 547774 153414 548354 188858
rect 547774 153178 547946 153414
rect 548182 153178 548354 153414
rect 547774 153094 548354 153178
rect 547774 152858 547946 153094
rect 548182 152858 548354 153094
rect 547774 117414 548354 152858
rect 547774 117178 547946 117414
rect 548182 117178 548354 117414
rect 547774 117094 548354 117178
rect 547774 116858 547946 117094
rect 548182 116858 548354 117094
rect 547774 81414 548354 116858
rect 547774 81178 547946 81414
rect 548182 81178 548354 81414
rect 547774 81094 548354 81178
rect 547774 80858 547946 81094
rect 548182 80858 548354 81094
rect 547774 45414 548354 80858
rect 547774 45178 547946 45414
rect 548182 45178 548354 45414
rect 547774 45094 548354 45178
rect 547774 44858 547946 45094
rect 548182 44858 548354 45094
rect 547774 9414 548354 44858
rect 547774 9178 547946 9414
rect 548182 9178 548354 9414
rect 547774 9094 548354 9178
rect 547774 8858 547946 9094
rect 548182 8858 548354 9094
rect 547774 -4026 548354 8858
rect 547774 -4262 547946 -4026
rect 548182 -4262 548354 -4026
rect 547774 -4346 548354 -4262
rect 547774 -4582 547946 -4346
rect 548182 -4582 548354 -4346
rect 547774 -5514 548354 -4582
rect 551254 696894 551834 709802
rect 569254 711278 569834 711290
rect 569254 711042 569426 711278
rect 569662 711042 569834 711278
rect 569254 710958 569834 711042
rect 569254 710722 569426 710958
rect 569662 710722 569834 710958
rect 565774 709438 566354 709450
rect 565774 709202 565946 709438
rect 566182 709202 566354 709438
rect 565774 709118 566354 709202
rect 565774 708882 565946 709118
rect 566182 708882 566354 709118
rect 562294 707598 562874 707610
rect 562294 707362 562466 707598
rect 562702 707362 562874 707598
rect 562294 707278 562874 707362
rect 562294 707042 562466 707278
rect 562702 707042 562874 707278
rect 551254 696658 551426 696894
rect 551662 696658 551834 696894
rect 551254 696574 551834 696658
rect 551254 696338 551426 696574
rect 551662 696338 551834 696574
rect 551254 660894 551834 696338
rect 551254 660658 551426 660894
rect 551662 660658 551834 660894
rect 551254 660574 551834 660658
rect 551254 660338 551426 660574
rect 551662 660338 551834 660574
rect 551254 624894 551834 660338
rect 551254 624658 551426 624894
rect 551662 624658 551834 624894
rect 551254 624574 551834 624658
rect 551254 624338 551426 624574
rect 551662 624338 551834 624574
rect 551254 588894 551834 624338
rect 551254 588658 551426 588894
rect 551662 588658 551834 588894
rect 551254 588574 551834 588658
rect 551254 588338 551426 588574
rect 551662 588338 551834 588574
rect 551254 552894 551834 588338
rect 551254 552658 551426 552894
rect 551662 552658 551834 552894
rect 551254 552574 551834 552658
rect 551254 552338 551426 552574
rect 551662 552338 551834 552574
rect 551254 516894 551834 552338
rect 551254 516658 551426 516894
rect 551662 516658 551834 516894
rect 551254 516574 551834 516658
rect 551254 516338 551426 516574
rect 551662 516338 551834 516574
rect 551254 480894 551834 516338
rect 551254 480658 551426 480894
rect 551662 480658 551834 480894
rect 551254 480574 551834 480658
rect 551254 480338 551426 480574
rect 551662 480338 551834 480574
rect 551254 444894 551834 480338
rect 551254 444658 551426 444894
rect 551662 444658 551834 444894
rect 551254 444574 551834 444658
rect 551254 444338 551426 444574
rect 551662 444338 551834 444574
rect 551254 408894 551834 444338
rect 551254 408658 551426 408894
rect 551662 408658 551834 408894
rect 551254 408574 551834 408658
rect 551254 408338 551426 408574
rect 551662 408338 551834 408574
rect 551254 372894 551834 408338
rect 551254 372658 551426 372894
rect 551662 372658 551834 372894
rect 551254 372574 551834 372658
rect 551254 372338 551426 372574
rect 551662 372338 551834 372574
rect 551254 336894 551834 372338
rect 551254 336658 551426 336894
rect 551662 336658 551834 336894
rect 551254 336574 551834 336658
rect 551254 336338 551426 336574
rect 551662 336338 551834 336574
rect 551254 300894 551834 336338
rect 551254 300658 551426 300894
rect 551662 300658 551834 300894
rect 551254 300574 551834 300658
rect 551254 300338 551426 300574
rect 551662 300338 551834 300574
rect 551254 264894 551834 300338
rect 551254 264658 551426 264894
rect 551662 264658 551834 264894
rect 551254 264574 551834 264658
rect 551254 264338 551426 264574
rect 551662 264338 551834 264574
rect 551254 228894 551834 264338
rect 551254 228658 551426 228894
rect 551662 228658 551834 228894
rect 551254 228574 551834 228658
rect 551254 228338 551426 228574
rect 551662 228338 551834 228574
rect 551254 192894 551834 228338
rect 551254 192658 551426 192894
rect 551662 192658 551834 192894
rect 551254 192574 551834 192658
rect 551254 192338 551426 192574
rect 551662 192338 551834 192574
rect 551254 156894 551834 192338
rect 551254 156658 551426 156894
rect 551662 156658 551834 156894
rect 551254 156574 551834 156658
rect 551254 156338 551426 156574
rect 551662 156338 551834 156574
rect 551254 120894 551834 156338
rect 551254 120658 551426 120894
rect 551662 120658 551834 120894
rect 551254 120574 551834 120658
rect 551254 120338 551426 120574
rect 551662 120338 551834 120574
rect 551254 84894 551834 120338
rect 551254 84658 551426 84894
rect 551662 84658 551834 84894
rect 551254 84574 551834 84658
rect 551254 84338 551426 84574
rect 551662 84338 551834 84574
rect 551254 48894 551834 84338
rect 551254 48658 551426 48894
rect 551662 48658 551834 48894
rect 551254 48574 551834 48658
rect 551254 48338 551426 48574
rect 551662 48338 551834 48574
rect 551254 12894 551834 48338
rect 551254 12658 551426 12894
rect 551662 12658 551834 12894
rect 551254 12574 551834 12658
rect 551254 12338 551426 12574
rect 551662 12338 551834 12574
rect 533254 -7022 533426 -6786
rect 533662 -7022 533834 -6786
rect 533254 -7106 533834 -7022
rect 533254 -7342 533426 -7106
rect 533662 -7342 533834 -7106
rect 533254 -7354 533834 -7342
rect 551254 -5866 551834 12338
rect 558814 705758 559394 705770
rect 558814 705522 558986 705758
rect 559222 705522 559394 705758
rect 558814 705438 559394 705522
rect 558814 705202 558986 705438
rect 559222 705202 559394 705438
rect 558814 668454 559394 705202
rect 558814 668218 558986 668454
rect 559222 668218 559394 668454
rect 558814 668134 559394 668218
rect 558814 667898 558986 668134
rect 559222 667898 559394 668134
rect 558814 632454 559394 667898
rect 558814 632218 558986 632454
rect 559222 632218 559394 632454
rect 558814 632134 559394 632218
rect 558814 631898 558986 632134
rect 559222 631898 559394 632134
rect 558814 596454 559394 631898
rect 558814 596218 558986 596454
rect 559222 596218 559394 596454
rect 558814 596134 559394 596218
rect 558814 595898 558986 596134
rect 559222 595898 559394 596134
rect 558814 560454 559394 595898
rect 558814 560218 558986 560454
rect 559222 560218 559394 560454
rect 558814 560134 559394 560218
rect 558814 559898 558986 560134
rect 559222 559898 559394 560134
rect 558814 524454 559394 559898
rect 558814 524218 558986 524454
rect 559222 524218 559394 524454
rect 558814 524134 559394 524218
rect 558814 523898 558986 524134
rect 559222 523898 559394 524134
rect 558814 488454 559394 523898
rect 558814 488218 558986 488454
rect 559222 488218 559394 488454
rect 558814 488134 559394 488218
rect 558814 487898 558986 488134
rect 559222 487898 559394 488134
rect 558814 452454 559394 487898
rect 558814 452218 558986 452454
rect 559222 452218 559394 452454
rect 558814 452134 559394 452218
rect 558814 451898 558986 452134
rect 559222 451898 559394 452134
rect 558814 416454 559394 451898
rect 558814 416218 558986 416454
rect 559222 416218 559394 416454
rect 558814 416134 559394 416218
rect 558814 415898 558986 416134
rect 559222 415898 559394 416134
rect 558814 380454 559394 415898
rect 558814 380218 558986 380454
rect 559222 380218 559394 380454
rect 558814 380134 559394 380218
rect 558814 379898 558986 380134
rect 559222 379898 559394 380134
rect 558814 344454 559394 379898
rect 558814 344218 558986 344454
rect 559222 344218 559394 344454
rect 558814 344134 559394 344218
rect 558814 343898 558986 344134
rect 559222 343898 559394 344134
rect 558814 308454 559394 343898
rect 558814 308218 558986 308454
rect 559222 308218 559394 308454
rect 558814 308134 559394 308218
rect 558814 307898 558986 308134
rect 559222 307898 559394 308134
rect 558814 272454 559394 307898
rect 558814 272218 558986 272454
rect 559222 272218 559394 272454
rect 558814 272134 559394 272218
rect 558814 271898 558986 272134
rect 559222 271898 559394 272134
rect 558814 236454 559394 271898
rect 558814 236218 558986 236454
rect 559222 236218 559394 236454
rect 558814 236134 559394 236218
rect 558814 235898 558986 236134
rect 559222 235898 559394 236134
rect 558814 200454 559394 235898
rect 558814 200218 558986 200454
rect 559222 200218 559394 200454
rect 558814 200134 559394 200218
rect 558814 199898 558986 200134
rect 559222 199898 559394 200134
rect 558814 164454 559394 199898
rect 558814 164218 558986 164454
rect 559222 164218 559394 164454
rect 558814 164134 559394 164218
rect 558814 163898 558986 164134
rect 559222 163898 559394 164134
rect 558814 128454 559394 163898
rect 558814 128218 558986 128454
rect 559222 128218 559394 128454
rect 558814 128134 559394 128218
rect 558814 127898 558986 128134
rect 559222 127898 559394 128134
rect 558814 92454 559394 127898
rect 558814 92218 558986 92454
rect 559222 92218 559394 92454
rect 558814 92134 559394 92218
rect 558814 91898 558986 92134
rect 559222 91898 559394 92134
rect 558814 56454 559394 91898
rect 558814 56218 558986 56454
rect 559222 56218 559394 56454
rect 558814 56134 559394 56218
rect 558814 55898 558986 56134
rect 559222 55898 559394 56134
rect 558814 20454 559394 55898
rect 558814 20218 558986 20454
rect 559222 20218 559394 20454
rect 558814 20134 559394 20218
rect 558814 19898 558986 20134
rect 559222 19898 559394 20134
rect 558814 -1266 559394 19898
rect 558814 -1502 558986 -1266
rect 559222 -1502 559394 -1266
rect 558814 -1586 559394 -1502
rect 558814 -1822 558986 -1586
rect 559222 -1822 559394 -1586
rect 558814 -1834 559394 -1822
rect 562294 671934 562874 707042
rect 562294 671698 562466 671934
rect 562702 671698 562874 671934
rect 562294 671614 562874 671698
rect 562294 671378 562466 671614
rect 562702 671378 562874 671614
rect 562294 635934 562874 671378
rect 562294 635698 562466 635934
rect 562702 635698 562874 635934
rect 562294 635614 562874 635698
rect 562294 635378 562466 635614
rect 562702 635378 562874 635614
rect 562294 599934 562874 635378
rect 562294 599698 562466 599934
rect 562702 599698 562874 599934
rect 562294 599614 562874 599698
rect 562294 599378 562466 599614
rect 562702 599378 562874 599614
rect 562294 563934 562874 599378
rect 562294 563698 562466 563934
rect 562702 563698 562874 563934
rect 562294 563614 562874 563698
rect 562294 563378 562466 563614
rect 562702 563378 562874 563614
rect 562294 527934 562874 563378
rect 562294 527698 562466 527934
rect 562702 527698 562874 527934
rect 562294 527614 562874 527698
rect 562294 527378 562466 527614
rect 562702 527378 562874 527614
rect 562294 491934 562874 527378
rect 562294 491698 562466 491934
rect 562702 491698 562874 491934
rect 562294 491614 562874 491698
rect 562294 491378 562466 491614
rect 562702 491378 562874 491614
rect 562294 455934 562874 491378
rect 562294 455698 562466 455934
rect 562702 455698 562874 455934
rect 562294 455614 562874 455698
rect 562294 455378 562466 455614
rect 562702 455378 562874 455614
rect 562294 419934 562874 455378
rect 562294 419698 562466 419934
rect 562702 419698 562874 419934
rect 562294 419614 562874 419698
rect 562294 419378 562466 419614
rect 562702 419378 562874 419614
rect 562294 383934 562874 419378
rect 562294 383698 562466 383934
rect 562702 383698 562874 383934
rect 562294 383614 562874 383698
rect 562294 383378 562466 383614
rect 562702 383378 562874 383614
rect 562294 347934 562874 383378
rect 562294 347698 562466 347934
rect 562702 347698 562874 347934
rect 562294 347614 562874 347698
rect 562294 347378 562466 347614
rect 562702 347378 562874 347614
rect 562294 311934 562874 347378
rect 562294 311698 562466 311934
rect 562702 311698 562874 311934
rect 562294 311614 562874 311698
rect 562294 311378 562466 311614
rect 562702 311378 562874 311614
rect 562294 275934 562874 311378
rect 562294 275698 562466 275934
rect 562702 275698 562874 275934
rect 562294 275614 562874 275698
rect 562294 275378 562466 275614
rect 562702 275378 562874 275614
rect 562294 239934 562874 275378
rect 562294 239698 562466 239934
rect 562702 239698 562874 239934
rect 562294 239614 562874 239698
rect 562294 239378 562466 239614
rect 562702 239378 562874 239614
rect 562294 203934 562874 239378
rect 562294 203698 562466 203934
rect 562702 203698 562874 203934
rect 562294 203614 562874 203698
rect 562294 203378 562466 203614
rect 562702 203378 562874 203614
rect 562294 167934 562874 203378
rect 562294 167698 562466 167934
rect 562702 167698 562874 167934
rect 562294 167614 562874 167698
rect 562294 167378 562466 167614
rect 562702 167378 562874 167614
rect 562294 131934 562874 167378
rect 562294 131698 562466 131934
rect 562702 131698 562874 131934
rect 562294 131614 562874 131698
rect 562294 131378 562466 131614
rect 562702 131378 562874 131614
rect 562294 95934 562874 131378
rect 562294 95698 562466 95934
rect 562702 95698 562874 95934
rect 562294 95614 562874 95698
rect 562294 95378 562466 95614
rect 562702 95378 562874 95614
rect 562294 59934 562874 95378
rect 562294 59698 562466 59934
rect 562702 59698 562874 59934
rect 562294 59614 562874 59698
rect 562294 59378 562466 59614
rect 562702 59378 562874 59614
rect 562294 23934 562874 59378
rect 562294 23698 562466 23934
rect 562702 23698 562874 23934
rect 562294 23614 562874 23698
rect 562294 23378 562466 23614
rect 562702 23378 562874 23614
rect 562294 -3106 562874 23378
rect 562294 -3342 562466 -3106
rect 562702 -3342 562874 -3106
rect 562294 -3426 562874 -3342
rect 562294 -3662 562466 -3426
rect 562702 -3662 562874 -3426
rect 562294 -3674 562874 -3662
rect 565774 675414 566354 708882
rect 565774 675178 565946 675414
rect 566182 675178 566354 675414
rect 565774 675094 566354 675178
rect 565774 674858 565946 675094
rect 566182 674858 566354 675094
rect 565774 639414 566354 674858
rect 565774 639178 565946 639414
rect 566182 639178 566354 639414
rect 565774 639094 566354 639178
rect 565774 638858 565946 639094
rect 566182 638858 566354 639094
rect 565774 603414 566354 638858
rect 565774 603178 565946 603414
rect 566182 603178 566354 603414
rect 565774 603094 566354 603178
rect 565774 602858 565946 603094
rect 566182 602858 566354 603094
rect 565774 567414 566354 602858
rect 565774 567178 565946 567414
rect 566182 567178 566354 567414
rect 565774 567094 566354 567178
rect 565774 566858 565946 567094
rect 566182 566858 566354 567094
rect 565774 531414 566354 566858
rect 565774 531178 565946 531414
rect 566182 531178 566354 531414
rect 565774 531094 566354 531178
rect 565774 530858 565946 531094
rect 566182 530858 566354 531094
rect 565774 495414 566354 530858
rect 565774 495178 565946 495414
rect 566182 495178 566354 495414
rect 565774 495094 566354 495178
rect 565774 494858 565946 495094
rect 566182 494858 566354 495094
rect 565774 459414 566354 494858
rect 565774 459178 565946 459414
rect 566182 459178 566354 459414
rect 565774 459094 566354 459178
rect 565774 458858 565946 459094
rect 566182 458858 566354 459094
rect 565774 423414 566354 458858
rect 565774 423178 565946 423414
rect 566182 423178 566354 423414
rect 565774 423094 566354 423178
rect 565774 422858 565946 423094
rect 566182 422858 566354 423094
rect 565774 387414 566354 422858
rect 565774 387178 565946 387414
rect 566182 387178 566354 387414
rect 565774 387094 566354 387178
rect 565774 386858 565946 387094
rect 566182 386858 566354 387094
rect 565774 351414 566354 386858
rect 565774 351178 565946 351414
rect 566182 351178 566354 351414
rect 565774 351094 566354 351178
rect 565774 350858 565946 351094
rect 566182 350858 566354 351094
rect 565774 315414 566354 350858
rect 565774 315178 565946 315414
rect 566182 315178 566354 315414
rect 565774 315094 566354 315178
rect 565774 314858 565946 315094
rect 566182 314858 566354 315094
rect 565774 279414 566354 314858
rect 565774 279178 565946 279414
rect 566182 279178 566354 279414
rect 565774 279094 566354 279178
rect 565774 278858 565946 279094
rect 566182 278858 566354 279094
rect 565774 243414 566354 278858
rect 565774 243178 565946 243414
rect 566182 243178 566354 243414
rect 565774 243094 566354 243178
rect 565774 242858 565946 243094
rect 566182 242858 566354 243094
rect 565774 207414 566354 242858
rect 565774 207178 565946 207414
rect 566182 207178 566354 207414
rect 565774 207094 566354 207178
rect 565774 206858 565946 207094
rect 566182 206858 566354 207094
rect 565774 171414 566354 206858
rect 565774 171178 565946 171414
rect 566182 171178 566354 171414
rect 565774 171094 566354 171178
rect 565774 170858 565946 171094
rect 566182 170858 566354 171094
rect 565774 135414 566354 170858
rect 565774 135178 565946 135414
rect 566182 135178 566354 135414
rect 565774 135094 566354 135178
rect 565774 134858 565946 135094
rect 566182 134858 566354 135094
rect 565774 99414 566354 134858
rect 565774 99178 565946 99414
rect 566182 99178 566354 99414
rect 565774 99094 566354 99178
rect 565774 98858 565946 99094
rect 566182 98858 566354 99094
rect 565774 63414 566354 98858
rect 565774 63178 565946 63414
rect 566182 63178 566354 63414
rect 565774 63094 566354 63178
rect 565774 62858 565946 63094
rect 566182 62858 566354 63094
rect 565774 27414 566354 62858
rect 565774 27178 565946 27414
rect 566182 27178 566354 27414
rect 565774 27094 566354 27178
rect 565774 26858 565946 27094
rect 566182 26858 566354 27094
rect 565774 -4946 566354 26858
rect 565774 -5182 565946 -4946
rect 566182 -5182 566354 -4946
rect 565774 -5266 566354 -5182
rect 565774 -5502 565946 -5266
rect 566182 -5502 566354 -5266
rect 565774 -5514 566354 -5502
rect 569254 678894 569834 710722
rect 591770 711278 592350 711290
rect 591770 711042 591942 711278
rect 592178 711042 592350 711278
rect 591770 710958 592350 711042
rect 591770 710722 591942 710958
rect 592178 710722 592350 710958
rect 590850 710358 591430 710370
rect 590850 710122 591022 710358
rect 591258 710122 591430 710358
rect 590850 710038 591430 710122
rect 590850 709802 591022 710038
rect 591258 709802 591430 710038
rect 589930 709438 590510 709450
rect 589930 709202 590102 709438
rect 590338 709202 590510 709438
rect 589930 709118 590510 709202
rect 589930 708882 590102 709118
rect 590338 708882 590510 709118
rect 589010 708518 589590 708530
rect 589010 708282 589182 708518
rect 589418 708282 589590 708518
rect 589010 708198 589590 708282
rect 589010 707962 589182 708198
rect 589418 707962 589590 708198
rect 580294 706678 580874 707610
rect 588090 707598 588670 707610
rect 588090 707362 588262 707598
rect 588498 707362 588670 707598
rect 588090 707278 588670 707362
rect 588090 707042 588262 707278
rect 588498 707042 588670 707278
rect 580294 706442 580466 706678
rect 580702 706442 580874 706678
rect 580294 706358 580874 706442
rect 580294 706122 580466 706358
rect 580702 706122 580874 706358
rect 569254 678658 569426 678894
rect 569662 678658 569834 678894
rect 569254 678574 569834 678658
rect 569254 678338 569426 678574
rect 569662 678338 569834 678574
rect 569254 642894 569834 678338
rect 569254 642658 569426 642894
rect 569662 642658 569834 642894
rect 569254 642574 569834 642658
rect 569254 642338 569426 642574
rect 569662 642338 569834 642574
rect 569254 606894 569834 642338
rect 569254 606658 569426 606894
rect 569662 606658 569834 606894
rect 569254 606574 569834 606658
rect 569254 606338 569426 606574
rect 569662 606338 569834 606574
rect 569254 570894 569834 606338
rect 569254 570658 569426 570894
rect 569662 570658 569834 570894
rect 569254 570574 569834 570658
rect 569254 570338 569426 570574
rect 569662 570338 569834 570574
rect 569254 534894 569834 570338
rect 569254 534658 569426 534894
rect 569662 534658 569834 534894
rect 569254 534574 569834 534658
rect 569254 534338 569426 534574
rect 569662 534338 569834 534574
rect 569254 498894 569834 534338
rect 569254 498658 569426 498894
rect 569662 498658 569834 498894
rect 569254 498574 569834 498658
rect 569254 498338 569426 498574
rect 569662 498338 569834 498574
rect 569254 462894 569834 498338
rect 569254 462658 569426 462894
rect 569662 462658 569834 462894
rect 569254 462574 569834 462658
rect 569254 462338 569426 462574
rect 569662 462338 569834 462574
rect 569254 426894 569834 462338
rect 569254 426658 569426 426894
rect 569662 426658 569834 426894
rect 569254 426574 569834 426658
rect 569254 426338 569426 426574
rect 569662 426338 569834 426574
rect 569254 390894 569834 426338
rect 569254 390658 569426 390894
rect 569662 390658 569834 390894
rect 569254 390574 569834 390658
rect 569254 390338 569426 390574
rect 569662 390338 569834 390574
rect 569254 354894 569834 390338
rect 569254 354658 569426 354894
rect 569662 354658 569834 354894
rect 569254 354574 569834 354658
rect 569254 354338 569426 354574
rect 569662 354338 569834 354574
rect 569254 318894 569834 354338
rect 569254 318658 569426 318894
rect 569662 318658 569834 318894
rect 569254 318574 569834 318658
rect 569254 318338 569426 318574
rect 569662 318338 569834 318574
rect 569254 282894 569834 318338
rect 569254 282658 569426 282894
rect 569662 282658 569834 282894
rect 569254 282574 569834 282658
rect 569254 282338 569426 282574
rect 569662 282338 569834 282574
rect 569254 246894 569834 282338
rect 569254 246658 569426 246894
rect 569662 246658 569834 246894
rect 569254 246574 569834 246658
rect 569254 246338 569426 246574
rect 569662 246338 569834 246574
rect 569254 210894 569834 246338
rect 569254 210658 569426 210894
rect 569662 210658 569834 210894
rect 569254 210574 569834 210658
rect 569254 210338 569426 210574
rect 569662 210338 569834 210574
rect 569254 174894 569834 210338
rect 569254 174658 569426 174894
rect 569662 174658 569834 174894
rect 569254 174574 569834 174658
rect 569254 174338 569426 174574
rect 569662 174338 569834 174574
rect 569254 138894 569834 174338
rect 569254 138658 569426 138894
rect 569662 138658 569834 138894
rect 569254 138574 569834 138658
rect 569254 138338 569426 138574
rect 569662 138338 569834 138574
rect 569254 102894 569834 138338
rect 569254 102658 569426 102894
rect 569662 102658 569834 102894
rect 569254 102574 569834 102658
rect 569254 102338 569426 102574
rect 569662 102338 569834 102574
rect 569254 66894 569834 102338
rect 569254 66658 569426 66894
rect 569662 66658 569834 66894
rect 569254 66574 569834 66658
rect 569254 66338 569426 66574
rect 569662 66338 569834 66574
rect 569254 30894 569834 66338
rect 569254 30658 569426 30894
rect 569662 30658 569834 30894
rect 569254 30574 569834 30658
rect 569254 30338 569426 30574
rect 569662 30338 569834 30574
rect 551254 -6102 551426 -5866
rect 551662 -6102 551834 -5866
rect 551254 -6186 551834 -6102
rect 551254 -6422 551426 -6186
rect 551662 -6422 551834 -6186
rect 551254 -7354 551834 -6422
rect 569254 -6786 569834 30338
rect 576814 704838 577394 705770
rect 576814 704602 576986 704838
rect 577222 704602 577394 704838
rect 576814 704518 577394 704602
rect 576814 704282 576986 704518
rect 577222 704282 577394 704518
rect 576814 686454 577394 704282
rect 576814 686218 576986 686454
rect 577222 686218 577394 686454
rect 576814 686134 577394 686218
rect 576814 685898 576986 686134
rect 577222 685898 577394 686134
rect 576814 650454 577394 685898
rect 576814 650218 576986 650454
rect 577222 650218 577394 650454
rect 576814 650134 577394 650218
rect 576814 649898 576986 650134
rect 577222 649898 577394 650134
rect 576814 614454 577394 649898
rect 576814 614218 576986 614454
rect 577222 614218 577394 614454
rect 576814 614134 577394 614218
rect 576814 613898 576986 614134
rect 577222 613898 577394 614134
rect 576814 578454 577394 613898
rect 576814 578218 576986 578454
rect 577222 578218 577394 578454
rect 576814 578134 577394 578218
rect 576814 577898 576986 578134
rect 577222 577898 577394 578134
rect 576814 542454 577394 577898
rect 576814 542218 576986 542454
rect 577222 542218 577394 542454
rect 576814 542134 577394 542218
rect 576814 541898 576986 542134
rect 577222 541898 577394 542134
rect 576814 506454 577394 541898
rect 576814 506218 576986 506454
rect 577222 506218 577394 506454
rect 576814 506134 577394 506218
rect 576814 505898 576986 506134
rect 577222 505898 577394 506134
rect 576814 470454 577394 505898
rect 576814 470218 576986 470454
rect 577222 470218 577394 470454
rect 576814 470134 577394 470218
rect 576814 469898 576986 470134
rect 577222 469898 577394 470134
rect 576814 434454 577394 469898
rect 576814 434218 576986 434454
rect 577222 434218 577394 434454
rect 576814 434134 577394 434218
rect 576814 433898 576986 434134
rect 577222 433898 577394 434134
rect 576814 398454 577394 433898
rect 576814 398218 576986 398454
rect 577222 398218 577394 398454
rect 576814 398134 577394 398218
rect 576814 397898 576986 398134
rect 577222 397898 577394 398134
rect 576814 362454 577394 397898
rect 576814 362218 576986 362454
rect 577222 362218 577394 362454
rect 576814 362134 577394 362218
rect 576814 361898 576986 362134
rect 577222 361898 577394 362134
rect 576814 326454 577394 361898
rect 576814 326218 576986 326454
rect 577222 326218 577394 326454
rect 576814 326134 577394 326218
rect 576814 325898 576986 326134
rect 577222 325898 577394 326134
rect 576814 290454 577394 325898
rect 576814 290218 576986 290454
rect 577222 290218 577394 290454
rect 576814 290134 577394 290218
rect 576814 289898 576986 290134
rect 577222 289898 577394 290134
rect 576814 254454 577394 289898
rect 576814 254218 576986 254454
rect 577222 254218 577394 254454
rect 576814 254134 577394 254218
rect 576814 253898 576986 254134
rect 577222 253898 577394 254134
rect 576814 218454 577394 253898
rect 576814 218218 576986 218454
rect 577222 218218 577394 218454
rect 576814 218134 577394 218218
rect 576814 217898 576986 218134
rect 577222 217898 577394 218134
rect 576814 182454 577394 217898
rect 576814 182218 576986 182454
rect 577222 182218 577394 182454
rect 576814 182134 577394 182218
rect 576814 181898 576986 182134
rect 577222 181898 577394 182134
rect 576814 146454 577394 181898
rect 576814 146218 576986 146454
rect 577222 146218 577394 146454
rect 576814 146134 577394 146218
rect 576814 145898 576986 146134
rect 577222 145898 577394 146134
rect 576814 110454 577394 145898
rect 576814 110218 576986 110454
rect 577222 110218 577394 110454
rect 576814 110134 577394 110218
rect 576814 109898 576986 110134
rect 577222 109898 577394 110134
rect 576814 74454 577394 109898
rect 576814 74218 576986 74454
rect 577222 74218 577394 74454
rect 576814 74134 577394 74218
rect 576814 73898 576986 74134
rect 577222 73898 577394 74134
rect 576814 38454 577394 73898
rect 576814 38218 576986 38454
rect 577222 38218 577394 38454
rect 576814 38134 577394 38218
rect 576814 37898 576986 38134
rect 577222 37898 577394 38134
rect 576814 2454 577394 37898
rect 576814 2218 576986 2454
rect 577222 2218 577394 2454
rect 576814 2134 577394 2218
rect 576814 1898 576986 2134
rect 577222 1898 577394 2134
rect 576814 -346 577394 1898
rect 576814 -582 576986 -346
rect 577222 -582 577394 -346
rect 576814 -666 577394 -582
rect 576814 -902 576986 -666
rect 577222 -902 577394 -666
rect 576814 -1834 577394 -902
rect 580294 689934 580874 706122
rect 587170 706678 587750 706690
rect 587170 706442 587342 706678
rect 587578 706442 587750 706678
rect 587170 706358 587750 706442
rect 587170 706122 587342 706358
rect 587578 706122 587750 706358
rect 586250 705758 586830 705770
rect 586250 705522 586422 705758
rect 586658 705522 586830 705758
rect 586250 705438 586830 705522
rect 586250 705202 586422 705438
rect 586658 705202 586830 705438
rect 580294 689698 580466 689934
rect 580702 689698 580874 689934
rect 580294 689614 580874 689698
rect 580294 689378 580466 689614
rect 580702 689378 580874 689614
rect 580294 653934 580874 689378
rect 580294 653698 580466 653934
rect 580702 653698 580874 653934
rect 580294 653614 580874 653698
rect 580294 653378 580466 653614
rect 580702 653378 580874 653614
rect 580294 617934 580874 653378
rect 580294 617698 580466 617934
rect 580702 617698 580874 617934
rect 580294 617614 580874 617698
rect 580294 617378 580466 617614
rect 580702 617378 580874 617614
rect 580294 581934 580874 617378
rect 580294 581698 580466 581934
rect 580702 581698 580874 581934
rect 580294 581614 580874 581698
rect 580294 581378 580466 581614
rect 580702 581378 580874 581614
rect 580294 545934 580874 581378
rect 580294 545698 580466 545934
rect 580702 545698 580874 545934
rect 580294 545614 580874 545698
rect 580294 545378 580466 545614
rect 580702 545378 580874 545614
rect 580294 509934 580874 545378
rect 580294 509698 580466 509934
rect 580702 509698 580874 509934
rect 580294 509614 580874 509698
rect 580294 509378 580466 509614
rect 580702 509378 580874 509614
rect 580294 473934 580874 509378
rect 580294 473698 580466 473934
rect 580702 473698 580874 473934
rect 580294 473614 580874 473698
rect 580294 473378 580466 473614
rect 580702 473378 580874 473614
rect 580294 437934 580874 473378
rect 580294 437698 580466 437934
rect 580702 437698 580874 437934
rect 580294 437614 580874 437698
rect 580294 437378 580466 437614
rect 580702 437378 580874 437614
rect 580294 401934 580874 437378
rect 580294 401698 580466 401934
rect 580702 401698 580874 401934
rect 580294 401614 580874 401698
rect 580294 401378 580466 401614
rect 580702 401378 580874 401614
rect 580294 365934 580874 401378
rect 580294 365698 580466 365934
rect 580702 365698 580874 365934
rect 580294 365614 580874 365698
rect 580294 365378 580466 365614
rect 580702 365378 580874 365614
rect 580294 329934 580874 365378
rect 580294 329698 580466 329934
rect 580702 329698 580874 329934
rect 580294 329614 580874 329698
rect 580294 329378 580466 329614
rect 580702 329378 580874 329614
rect 580294 293934 580874 329378
rect 580294 293698 580466 293934
rect 580702 293698 580874 293934
rect 580294 293614 580874 293698
rect 580294 293378 580466 293614
rect 580702 293378 580874 293614
rect 580294 257934 580874 293378
rect 580294 257698 580466 257934
rect 580702 257698 580874 257934
rect 580294 257614 580874 257698
rect 580294 257378 580466 257614
rect 580702 257378 580874 257614
rect 580294 221934 580874 257378
rect 580294 221698 580466 221934
rect 580702 221698 580874 221934
rect 580294 221614 580874 221698
rect 580294 221378 580466 221614
rect 580702 221378 580874 221614
rect 580294 185934 580874 221378
rect 580294 185698 580466 185934
rect 580702 185698 580874 185934
rect 580294 185614 580874 185698
rect 580294 185378 580466 185614
rect 580702 185378 580874 185614
rect 580294 149934 580874 185378
rect 580294 149698 580466 149934
rect 580702 149698 580874 149934
rect 580294 149614 580874 149698
rect 580294 149378 580466 149614
rect 580702 149378 580874 149614
rect 580294 113934 580874 149378
rect 580294 113698 580466 113934
rect 580702 113698 580874 113934
rect 580294 113614 580874 113698
rect 580294 113378 580466 113614
rect 580702 113378 580874 113614
rect 580294 77934 580874 113378
rect 580294 77698 580466 77934
rect 580702 77698 580874 77934
rect 580294 77614 580874 77698
rect 580294 77378 580466 77614
rect 580702 77378 580874 77614
rect 580294 41934 580874 77378
rect 580294 41698 580466 41934
rect 580702 41698 580874 41934
rect 580294 41614 580874 41698
rect 580294 41378 580466 41614
rect 580702 41378 580874 41614
rect 580294 5934 580874 41378
rect 580294 5698 580466 5934
rect 580702 5698 580874 5934
rect 580294 5614 580874 5698
rect 580294 5378 580466 5614
rect 580702 5378 580874 5614
rect 580294 -2186 580874 5378
rect 585330 704838 585910 704850
rect 585330 704602 585502 704838
rect 585738 704602 585910 704838
rect 585330 704518 585910 704602
rect 585330 704282 585502 704518
rect 585738 704282 585910 704518
rect 585330 686454 585910 704282
rect 585330 686218 585502 686454
rect 585738 686218 585910 686454
rect 585330 686134 585910 686218
rect 585330 685898 585502 686134
rect 585738 685898 585910 686134
rect 585330 650454 585910 685898
rect 585330 650218 585502 650454
rect 585738 650218 585910 650454
rect 585330 650134 585910 650218
rect 585330 649898 585502 650134
rect 585738 649898 585910 650134
rect 585330 614454 585910 649898
rect 585330 614218 585502 614454
rect 585738 614218 585910 614454
rect 585330 614134 585910 614218
rect 585330 613898 585502 614134
rect 585738 613898 585910 614134
rect 585330 578454 585910 613898
rect 585330 578218 585502 578454
rect 585738 578218 585910 578454
rect 585330 578134 585910 578218
rect 585330 577898 585502 578134
rect 585738 577898 585910 578134
rect 585330 542454 585910 577898
rect 585330 542218 585502 542454
rect 585738 542218 585910 542454
rect 585330 542134 585910 542218
rect 585330 541898 585502 542134
rect 585738 541898 585910 542134
rect 585330 506454 585910 541898
rect 585330 506218 585502 506454
rect 585738 506218 585910 506454
rect 585330 506134 585910 506218
rect 585330 505898 585502 506134
rect 585738 505898 585910 506134
rect 585330 470454 585910 505898
rect 585330 470218 585502 470454
rect 585738 470218 585910 470454
rect 585330 470134 585910 470218
rect 585330 469898 585502 470134
rect 585738 469898 585910 470134
rect 585330 434454 585910 469898
rect 585330 434218 585502 434454
rect 585738 434218 585910 434454
rect 585330 434134 585910 434218
rect 585330 433898 585502 434134
rect 585738 433898 585910 434134
rect 585330 398454 585910 433898
rect 585330 398218 585502 398454
rect 585738 398218 585910 398454
rect 585330 398134 585910 398218
rect 585330 397898 585502 398134
rect 585738 397898 585910 398134
rect 585330 362454 585910 397898
rect 585330 362218 585502 362454
rect 585738 362218 585910 362454
rect 585330 362134 585910 362218
rect 585330 361898 585502 362134
rect 585738 361898 585910 362134
rect 585330 326454 585910 361898
rect 585330 326218 585502 326454
rect 585738 326218 585910 326454
rect 585330 326134 585910 326218
rect 585330 325898 585502 326134
rect 585738 325898 585910 326134
rect 585330 290454 585910 325898
rect 585330 290218 585502 290454
rect 585738 290218 585910 290454
rect 585330 290134 585910 290218
rect 585330 289898 585502 290134
rect 585738 289898 585910 290134
rect 585330 254454 585910 289898
rect 585330 254218 585502 254454
rect 585738 254218 585910 254454
rect 585330 254134 585910 254218
rect 585330 253898 585502 254134
rect 585738 253898 585910 254134
rect 585330 218454 585910 253898
rect 585330 218218 585502 218454
rect 585738 218218 585910 218454
rect 585330 218134 585910 218218
rect 585330 217898 585502 218134
rect 585738 217898 585910 218134
rect 585330 182454 585910 217898
rect 585330 182218 585502 182454
rect 585738 182218 585910 182454
rect 585330 182134 585910 182218
rect 585330 181898 585502 182134
rect 585738 181898 585910 182134
rect 585330 146454 585910 181898
rect 585330 146218 585502 146454
rect 585738 146218 585910 146454
rect 585330 146134 585910 146218
rect 585330 145898 585502 146134
rect 585738 145898 585910 146134
rect 585330 110454 585910 145898
rect 585330 110218 585502 110454
rect 585738 110218 585910 110454
rect 585330 110134 585910 110218
rect 585330 109898 585502 110134
rect 585738 109898 585910 110134
rect 585330 74454 585910 109898
rect 585330 74218 585502 74454
rect 585738 74218 585910 74454
rect 585330 74134 585910 74218
rect 585330 73898 585502 74134
rect 585738 73898 585910 74134
rect 585330 38454 585910 73898
rect 585330 38218 585502 38454
rect 585738 38218 585910 38454
rect 585330 38134 585910 38218
rect 585330 37898 585502 38134
rect 585738 37898 585910 38134
rect 585330 2454 585910 37898
rect 585330 2218 585502 2454
rect 585738 2218 585910 2454
rect 585330 2134 585910 2218
rect 585330 1898 585502 2134
rect 585738 1898 585910 2134
rect 585330 -346 585910 1898
rect 585330 -582 585502 -346
rect 585738 -582 585910 -346
rect 585330 -666 585910 -582
rect 585330 -902 585502 -666
rect 585738 -902 585910 -666
rect 585330 -914 585910 -902
rect 586250 668454 586830 705202
rect 586250 668218 586422 668454
rect 586658 668218 586830 668454
rect 586250 668134 586830 668218
rect 586250 667898 586422 668134
rect 586658 667898 586830 668134
rect 586250 632454 586830 667898
rect 586250 632218 586422 632454
rect 586658 632218 586830 632454
rect 586250 632134 586830 632218
rect 586250 631898 586422 632134
rect 586658 631898 586830 632134
rect 586250 596454 586830 631898
rect 586250 596218 586422 596454
rect 586658 596218 586830 596454
rect 586250 596134 586830 596218
rect 586250 595898 586422 596134
rect 586658 595898 586830 596134
rect 586250 560454 586830 595898
rect 586250 560218 586422 560454
rect 586658 560218 586830 560454
rect 586250 560134 586830 560218
rect 586250 559898 586422 560134
rect 586658 559898 586830 560134
rect 586250 524454 586830 559898
rect 586250 524218 586422 524454
rect 586658 524218 586830 524454
rect 586250 524134 586830 524218
rect 586250 523898 586422 524134
rect 586658 523898 586830 524134
rect 586250 488454 586830 523898
rect 586250 488218 586422 488454
rect 586658 488218 586830 488454
rect 586250 488134 586830 488218
rect 586250 487898 586422 488134
rect 586658 487898 586830 488134
rect 586250 452454 586830 487898
rect 586250 452218 586422 452454
rect 586658 452218 586830 452454
rect 586250 452134 586830 452218
rect 586250 451898 586422 452134
rect 586658 451898 586830 452134
rect 586250 416454 586830 451898
rect 586250 416218 586422 416454
rect 586658 416218 586830 416454
rect 586250 416134 586830 416218
rect 586250 415898 586422 416134
rect 586658 415898 586830 416134
rect 586250 380454 586830 415898
rect 586250 380218 586422 380454
rect 586658 380218 586830 380454
rect 586250 380134 586830 380218
rect 586250 379898 586422 380134
rect 586658 379898 586830 380134
rect 586250 344454 586830 379898
rect 586250 344218 586422 344454
rect 586658 344218 586830 344454
rect 586250 344134 586830 344218
rect 586250 343898 586422 344134
rect 586658 343898 586830 344134
rect 586250 308454 586830 343898
rect 586250 308218 586422 308454
rect 586658 308218 586830 308454
rect 586250 308134 586830 308218
rect 586250 307898 586422 308134
rect 586658 307898 586830 308134
rect 586250 272454 586830 307898
rect 586250 272218 586422 272454
rect 586658 272218 586830 272454
rect 586250 272134 586830 272218
rect 586250 271898 586422 272134
rect 586658 271898 586830 272134
rect 586250 236454 586830 271898
rect 586250 236218 586422 236454
rect 586658 236218 586830 236454
rect 586250 236134 586830 236218
rect 586250 235898 586422 236134
rect 586658 235898 586830 236134
rect 586250 200454 586830 235898
rect 586250 200218 586422 200454
rect 586658 200218 586830 200454
rect 586250 200134 586830 200218
rect 586250 199898 586422 200134
rect 586658 199898 586830 200134
rect 586250 164454 586830 199898
rect 586250 164218 586422 164454
rect 586658 164218 586830 164454
rect 586250 164134 586830 164218
rect 586250 163898 586422 164134
rect 586658 163898 586830 164134
rect 586250 128454 586830 163898
rect 586250 128218 586422 128454
rect 586658 128218 586830 128454
rect 586250 128134 586830 128218
rect 586250 127898 586422 128134
rect 586658 127898 586830 128134
rect 586250 92454 586830 127898
rect 586250 92218 586422 92454
rect 586658 92218 586830 92454
rect 586250 92134 586830 92218
rect 586250 91898 586422 92134
rect 586658 91898 586830 92134
rect 586250 56454 586830 91898
rect 586250 56218 586422 56454
rect 586658 56218 586830 56454
rect 586250 56134 586830 56218
rect 586250 55898 586422 56134
rect 586658 55898 586830 56134
rect 586250 20454 586830 55898
rect 586250 20218 586422 20454
rect 586658 20218 586830 20454
rect 586250 20134 586830 20218
rect 586250 19898 586422 20134
rect 586658 19898 586830 20134
rect 586250 -1266 586830 19898
rect 586250 -1502 586422 -1266
rect 586658 -1502 586830 -1266
rect 586250 -1586 586830 -1502
rect 586250 -1822 586422 -1586
rect 586658 -1822 586830 -1586
rect 586250 -1834 586830 -1822
rect 587170 689934 587750 706122
rect 587170 689698 587342 689934
rect 587578 689698 587750 689934
rect 587170 689614 587750 689698
rect 587170 689378 587342 689614
rect 587578 689378 587750 689614
rect 587170 653934 587750 689378
rect 587170 653698 587342 653934
rect 587578 653698 587750 653934
rect 587170 653614 587750 653698
rect 587170 653378 587342 653614
rect 587578 653378 587750 653614
rect 587170 617934 587750 653378
rect 587170 617698 587342 617934
rect 587578 617698 587750 617934
rect 587170 617614 587750 617698
rect 587170 617378 587342 617614
rect 587578 617378 587750 617614
rect 587170 581934 587750 617378
rect 587170 581698 587342 581934
rect 587578 581698 587750 581934
rect 587170 581614 587750 581698
rect 587170 581378 587342 581614
rect 587578 581378 587750 581614
rect 587170 545934 587750 581378
rect 587170 545698 587342 545934
rect 587578 545698 587750 545934
rect 587170 545614 587750 545698
rect 587170 545378 587342 545614
rect 587578 545378 587750 545614
rect 587170 509934 587750 545378
rect 587170 509698 587342 509934
rect 587578 509698 587750 509934
rect 587170 509614 587750 509698
rect 587170 509378 587342 509614
rect 587578 509378 587750 509614
rect 587170 473934 587750 509378
rect 587170 473698 587342 473934
rect 587578 473698 587750 473934
rect 587170 473614 587750 473698
rect 587170 473378 587342 473614
rect 587578 473378 587750 473614
rect 587170 437934 587750 473378
rect 587170 437698 587342 437934
rect 587578 437698 587750 437934
rect 587170 437614 587750 437698
rect 587170 437378 587342 437614
rect 587578 437378 587750 437614
rect 587170 401934 587750 437378
rect 587170 401698 587342 401934
rect 587578 401698 587750 401934
rect 587170 401614 587750 401698
rect 587170 401378 587342 401614
rect 587578 401378 587750 401614
rect 587170 365934 587750 401378
rect 587170 365698 587342 365934
rect 587578 365698 587750 365934
rect 587170 365614 587750 365698
rect 587170 365378 587342 365614
rect 587578 365378 587750 365614
rect 587170 329934 587750 365378
rect 587170 329698 587342 329934
rect 587578 329698 587750 329934
rect 587170 329614 587750 329698
rect 587170 329378 587342 329614
rect 587578 329378 587750 329614
rect 587170 293934 587750 329378
rect 587170 293698 587342 293934
rect 587578 293698 587750 293934
rect 587170 293614 587750 293698
rect 587170 293378 587342 293614
rect 587578 293378 587750 293614
rect 587170 257934 587750 293378
rect 587170 257698 587342 257934
rect 587578 257698 587750 257934
rect 587170 257614 587750 257698
rect 587170 257378 587342 257614
rect 587578 257378 587750 257614
rect 587170 221934 587750 257378
rect 587170 221698 587342 221934
rect 587578 221698 587750 221934
rect 587170 221614 587750 221698
rect 587170 221378 587342 221614
rect 587578 221378 587750 221614
rect 587170 185934 587750 221378
rect 587170 185698 587342 185934
rect 587578 185698 587750 185934
rect 587170 185614 587750 185698
rect 587170 185378 587342 185614
rect 587578 185378 587750 185614
rect 587170 149934 587750 185378
rect 587170 149698 587342 149934
rect 587578 149698 587750 149934
rect 587170 149614 587750 149698
rect 587170 149378 587342 149614
rect 587578 149378 587750 149614
rect 587170 113934 587750 149378
rect 587170 113698 587342 113934
rect 587578 113698 587750 113934
rect 587170 113614 587750 113698
rect 587170 113378 587342 113614
rect 587578 113378 587750 113614
rect 587170 77934 587750 113378
rect 587170 77698 587342 77934
rect 587578 77698 587750 77934
rect 587170 77614 587750 77698
rect 587170 77378 587342 77614
rect 587578 77378 587750 77614
rect 587170 41934 587750 77378
rect 587170 41698 587342 41934
rect 587578 41698 587750 41934
rect 587170 41614 587750 41698
rect 587170 41378 587342 41614
rect 587578 41378 587750 41614
rect 587170 5934 587750 41378
rect 587170 5698 587342 5934
rect 587578 5698 587750 5934
rect 587170 5614 587750 5698
rect 587170 5378 587342 5614
rect 587578 5378 587750 5614
rect 580294 -2422 580466 -2186
rect 580702 -2422 580874 -2186
rect 580294 -2506 580874 -2422
rect 580294 -2742 580466 -2506
rect 580702 -2742 580874 -2506
rect 580294 -3674 580874 -2742
rect 587170 -2186 587750 5378
rect 587170 -2422 587342 -2186
rect 587578 -2422 587750 -2186
rect 587170 -2506 587750 -2422
rect 587170 -2742 587342 -2506
rect 587578 -2742 587750 -2506
rect 587170 -2754 587750 -2742
rect 588090 671934 588670 707042
rect 588090 671698 588262 671934
rect 588498 671698 588670 671934
rect 588090 671614 588670 671698
rect 588090 671378 588262 671614
rect 588498 671378 588670 671614
rect 588090 635934 588670 671378
rect 588090 635698 588262 635934
rect 588498 635698 588670 635934
rect 588090 635614 588670 635698
rect 588090 635378 588262 635614
rect 588498 635378 588670 635614
rect 588090 599934 588670 635378
rect 588090 599698 588262 599934
rect 588498 599698 588670 599934
rect 588090 599614 588670 599698
rect 588090 599378 588262 599614
rect 588498 599378 588670 599614
rect 588090 563934 588670 599378
rect 588090 563698 588262 563934
rect 588498 563698 588670 563934
rect 588090 563614 588670 563698
rect 588090 563378 588262 563614
rect 588498 563378 588670 563614
rect 588090 527934 588670 563378
rect 588090 527698 588262 527934
rect 588498 527698 588670 527934
rect 588090 527614 588670 527698
rect 588090 527378 588262 527614
rect 588498 527378 588670 527614
rect 588090 491934 588670 527378
rect 588090 491698 588262 491934
rect 588498 491698 588670 491934
rect 588090 491614 588670 491698
rect 588090 491378 588262 491614
rect 588498 491378 588670 491614
rect 588090 455934 588670 491378
rect 588090 455698 588262 455934
rect 588498 455698 588670 455934
rect 588090 455614 588670 455698
rect 588090 455378 588262 455614
rect 588498 455378 588670 455614
rect 588090 419934 588670 455378
rect 588090 419698 588262 419934
rect 588498 419698 588670 419934
rect 588090 419614 588670 419698
rect 588090 419378 588262 419614
rect 588498 419378 588670 419614
rect 588090 383934 588670 419378
rect 588090 383698 588262 383934
rect 588498 383698 588670 383934
rect 588090 383614 588670 383698
rect 588090 383378 588262 383614
rect 588498 383378 588670 383614
rect 588090 347934 588670 383378
rect 588090 347698 588262 347934
rect 588498 347698 588670 347934
rect 588090 347614 588670 347698
rect 588090 347378 588262 347614
rect 588498 347378 588670 347614
rect 588090 311934 588670 347378
rect 588090 311698 588262 311934
rect 588498 311698 588670 311934
rect 588090 311614 588670 311698
rect 588090 311378 588262 311614
rect 588498 311378 588670 311614
rect 588090 275934 588670 311378
rect 588090 275698 588262 275934
rect 588498 275698 588670 275934
rect 588090 275614 588670 275698
rect 588090 275378 588262 275614
rect 588498 275378 588670 275614
rect 588090 239934 588670 275378
rect 588090 239698 588262 239934
rect 588498 239698 588670 239934
rect 588090 239614 588670 239698
rect 588090 239378 588262 239614
rect 588498 239378 588670 239614
rect 588090 203934 588670 239378
rect 588090 203698 588262 203934
rect 588498 203698 588670 203934
rect 588090 203614 588670 203698
rect 588090 203378 588262 203614
rect 588498 203378 588670 203614
rect 588090 167934 588670 203378
rect 588090 167698 588262 167934
rect 588498 167698 588670 167934
rect 588090 167614 588670 167698
rect 588090 167378 588262 167614
rect 588498 167378 588670 167614
rect 588090 131934 588670 167378
rect 588090 131698 588262 131934
rect 588498 131698 588670 131934
rect 588090 131614 588670 131698
rect 588090 131378 588262 131614
rect 588498 131378 588670 131614
rect 588090 95934 588670 131378
rect 588090 95698 588262 95934
rect 588498 95698 588670 95934
rect 588090 95614 588670 95698
rect 588090 95378 588262 95614
rect 588498 95378 588670 95614
rect 588090 59934 588670 95378
rect 588090 59698 588262 59934
rect 588498 59698 588670 59934
rect 588090 59614 588670 59698
rect 588090 59378 588262 59614
rect 588498 59378 588670 59614
rect 588090 23934 588670 59378
rect 588090 23698 588262 23934
rect 588498 23698 588670 23934
rect 588090 23614 588670 23698
rect 588090 23378 588262 23614
rect 588498 23378 588670 23614
rect 588090 -3106 588670 23378
rect 588090 -3342 588262 -3106
rect 588498 -3342 588670 -3106
rect 588090 -3426 588670 -3342
rect 588090 -3662 588262 -3426
rect 588498 -3662 588670 -3426
rect 588090 -3674 588670 -3662
rect 589010 693414 589590 707962
rect 589010 693178 589182 693414
rect 589418 693178 589590 693414
rect 589010 693094 589590 693178
rect 589010 692858 589182 693094
rect 589418 692858 589590 693094
rect 589010 657414 589590 692858
rect 589010 657178 589182 657414
rect 589418 657178 589590 657414
rect 589010 657094 589590 657178
rect 589010 656858 589182 657094
rect 589418 656858 589590 657094
rect 589010 621414 589590 656858
rect 589010 621178 589182 621414
rect 589418 621178 589590 621414
rect 589010 621094 589590 621178
rect 589010 620858 589182 621094
rect 589418 620858 589590 621094
rect 589010 585414 589590 620858
rect 589010 585178 589182 585414
rect 589418 585178 589590 585414
rect 589010 585094 589590 585178
rect 589010 584858 589182 585094
rect 589418 584858 589590 585094
rect 589010 549414 589590 584858
rect 589010 549178 589182 549414
rect 589418 549178 589590 549414
rect 589010 549094 589590 549178
rect 589010 548858 589182 549094
rect 589418 548858 589590 549094
rect 589010 513414 589590 548858
rect 589010 513178 589182 513414
rect 589418 513178 589590 513414
rect 589010 513094 589590 513178
rect 589010 512858 589182 513094
rect 589418 512858 589590 513094
rect 589010 477414 589590 512858
rect 589010 477178 589182 477414
rect 589418 477178 589590 477414
rect 589010 477094 589590 477178
rect 589010 476858 589182 477094
rect 589418 476858 589590 477094
rect 589010 441414 589590 476858
rect 589010 441178 589182 441414
rect 589418 441178 589590 441414
rect 589010 441094 589590 441178
rect 589010 440858 589182 441094
rect 589418 440858 589590 441094
rect 589010 405414 589590 440858
rect 589010 405178 589182 405414
rect 589418 405178 589590 405414
rect 589010 405094 589590 405178
rect 589010 404858 589182 405094
rect 589418 404858 589590 405094
rect 589010 369414 589590 404858
rect 589010 369178 589182 369414
rect 589418 369178 589590 369414
rect 589010 369094 589590 369178
rect 589010 368858 589182 369094
rect 589418 368858 589590 369094
rect 589010 333414 589590 368858
rect 589010 333178 589182 333414
rect 589418 333178 589590 333414
rect 589010 333094 589590 333178
rect 589010 332858 589182 333094
rect 589418 332858 589590 333094
rect 589010 297414 589590 332858
rect 589010 297178 589182 297414
rect 589418 297178 589590 297414
rect 589010 297094 589590 297178
rect 589010 296858 589182 297094
rect 589418 296858 589590 297094
rect 589010 261414 589590 296858
rect 589010 261178 589182 261414
rect 589418 261178 589590 261414
rect 589010 261094 589590 261178
rect 589010 260858 589182 261094
rect 589418 260858 589590 261094
rect 589010 225414 589590 260858
rect 589010 225178 589182 225414
rect 589418 225178 589590 225414
rect 589010 225094 589590 225178
rect 589010 224858 589182 225094
rect 589418 224858 589590 225094
rect 589010 189414 589590 224858
rect 589010 189178 589182 189414
rect 589418 189178 589590 189414
rect 589010 189094 589590 189178
rect 589010 188858 589182 189094
rect 589418 188858 589590 189094
rect 589010 153414 589590 188858
rect 589010 153178 589182 153414
rect 589418 153178 589590 153414
rect 589010 153094 589590 153178
rect 589010 152858 589182 153094
rect 589418 152858 589590 153094
rect 589010 117414 589590 152858
rect 589010 117178 589182 117414
rect 589418 117178 589590 117414
rect 589010 117094 589590 117178
rect 589010 116858 589182 117094
rect 589418 116858 589590 117094
rect 589010 81414 589590 116858
rect 589010 81178 589182 81414
rect 589418 81178 589590 81414
rect 589010 81094 589590 81178
rect 589010 80858 589182 81094
rect 589418 80858 589590 81094
rect 589010 45414 589590 80858
rect 589010 45178 589182 45414
rect 589418 45178 589590 45414
rect 589010 45094 589590 45178
rect 589010 44858 589182 45094
rect 589418 44858 589590 45094
rect 589010 9414 589590 44858
rect 589010 9178 589182 9414
rect 589418 9178 589590 9414
rect 589010 9094 589590 9178
rect 589010 8858 589182 9094
rect 589418 8858 589590 9094
rect 589010 -4026 589590 8858
rect 589010 -4262 589182 -4026
rect 589418 -4262 589590 -4026
rect 589010 -4346 589590 -4262
rect 589010 -4582 589182 -4346
rect 589418 -4582 589590 -4346
rect 589010 -4594 589590 -4582
rect 589930 675414 590510 708882
rect 589930 675178 590102 675414
rect 590338 675178 590510 675414
rect 589930 675094 590510 675178
rect 589930 674858 590102 675094
rect 590338 674858 590510 675094
rect 589930 639414 590510 674858
rect 589930 639178 590102 639414
rect 590338 639178 590510 639414
rect 589930 639094 590510 639178
rect 589930 638858 590102 639094
rect 590338 638858 590510 639094
rect 589930 603414 590510 638858
rect 589930 603178 590102 603414
rect 590338 603178 590510 603414
rect 589930 603094 590510 603178
rect 589930 602858 590102 603094
rect 590338 602858 590510 603094
rect 589930 567414 590510 602858
rect 589930 567178 590102 567414
rect 590338 567178 590510 567414
rect 589930 567094 590510 567178
rect 589930 566858 590102 567094
rect 590338 566858 590510 567094
rect 589930 531414 590510 566858
rect 589930 531178 590102 531414
rect 590338 531178 590510 531414
rect 589930 531094 590510 531178
rect 589930 530858 590102 531094
rect 590338 530858 590510 531094
rect 589930 495414 590510 530858
rect 589930 495178 590102 495414
rect 590338 495178 590510 495414
rect 589930 495094 590510 495178
rect 589930 494858 590102 495094
rect 590338 494858 590510 495094
rect 589930 459414 590510 494858
rect 589930 459178 590102 459414
rect 590338 459178 590510 459414
rect 589930 459094 590510 459178
rect 589930 458858 590102 459094
rect 590338 458858 590510 459094
rect 589930 423414 590510 458858
rect 589930 423178 590102 423414
rect 590338 423178 590510 423414
rect 589930 423094 590510 423178
rect 589930 422858 590102 423094
rect 590338 422858 590510 423094
rect 589930 387414 590510 422858
rect 589930 387178 590102 387414
rect 590338 387178 590510 387414
rect 589930 387094 590510 387178
rect 589930 386858 590102 387094
rect 590338 386858 590510 387094
rect 589930 351414 590510 386858
rect 589930 351178 590102 351414
rect 590338 351178 590510 351414
rect 589930 351094 590510 351178
rect 589930 350858 590102 351094
rect 590338 350858 590510 351094
rect 589930 315414 590510 350858
rect 589930 315178 590102 315414
rect 590338 315178 590510 315414
rect 589930 315094 590510 315178
rect 589930 314858 590102 315094
rect 590338 314858 590510 315094
rect 589930 279414 590510 314858
rect 589930 279178 590102 279414
rect 590338 279178 590510 279414
rect 589930 279094 590510 279178
rect 589930 278858 590102 279094
rect 590338 278858 590510 279094
rect 589930 243414 590510 278858
rect 589930 243178 590102 243414
rect 590338 243178 590510 243414
rect 589930 243094 590510 243178
rect 589930 242858 590102 243094
rect 590338 242858 590510 243094
rect 589930 207414 590510 242858
rect 589930 207178 590102 207414
rect 590338 207178 590510 207414
rect 589930 207094 590510 207178
rect 589930 206858 590102 207094
rect 590338 206858 590510 207094
rect 589930 171414 590510 206858
rect 589930 171178 590102 171414
rect 590338 171178 590510 171414
rect 589930 171094 590510 171178
rect 589930 170858 590102 171094
rect 590338 170858 590510 171094
rect 589930 135414 590510 170858
rect 589930 135178 590102 135414
rect 590338 135178 590510 135414
rect 589930 135094 590510 135178
rect 589930 134858 590102 135094
rect 590338 134858 590510 135094
rect 589930 99414 590510 134858
rect 589930 99178 590102 99414
rect 590338 99178 590510 99414
rect 589930 99094 590510 99178
rect 589930 98858 590102 99094
rect 590338 98858 590510 99094
rect 589930 63414 590510 98858
rect 589930 63178 590102 63414
rect 590338 63178 590510 63414
rect 589930 63094 590510 63178
rect 589930 62858 590102 63094
rect 590338 62858 590510 63094
rect 589930 27414 590510 62858
rect 589930 27178 590102 27414
rect 590338 27178 590510 27414
rect 589930 27094 590510 27178
rect 589930 26858 590102 27094
rect 590338 26858 590510 27094
rect 589930 -4946 590510 26858
rect 589930 -5182 590102 -4946
rect 590338 -5182 590510 -4946
rect 589930 -5266 590510 -5182
rect 589930 -5502 590102 -5266
rect 590338 -5502 590510 -5266
rect 589930 -5514 590510 -5502
rect 590850 696894 591430 709802
rect 590850 696658 591022 696894
rect 591258 696658 591430 696894
rect 590850 696574 591430 696658
rect 590850 696338 591022 696574
rect 591258 696338 591430 696574
rect 590850 660894 591430 696338
rect 590850 660658 591022 660894
rect 591258 660658 591430 660894
rect 590850 660574 591430 660658
rect 590850 660338 591022 660574
rect 591258 660338 591430 660574
rect 590850 624894 591430 660338
rect 590850 624658 591022 624894
rect 591258 624658 591430 624894
rect 590850 624574 591430 624658
rect 590850 624338 591022 624574
rect 591258 624338 591430 624574
rect 590850 588894 591430 624338
rect 590850 588658 591022 588894
rect 591258 588658 591430 588894
rect 590850 588574 591430 588658
rect 590850 588338 591022 588574
rect 591258 588338 591430 588574
rect 590850 552894 591430 588338
rect 590850 552658 591022 552894
rect 591258 552658 591430 552894
rect 590850 552574 591430 552658
rect 590850 552338 591022 552574
rect 591258 552338 591430 552574
rect 590850 516894 591430 552338
rect 590850 516658 591022 516894
rect 591258 516658 591430 516894
rect 590850 516574 591430 516658
rect 590850 516338 591022 516574
rect 591258 516338 591430 516574
rect 590850 480894 591430 516338
rect 590850 480658 591022 480894
rect 591258 480658 591430 480894
rect 590850 480574 591430 480658
rect 590850 480338 591022 480574
rect 591258 480338 591430 480574
rect 590850 444894 591430 480338
rect 590850 444658 591022 444894
rect 591258 444658 591430 444894
rect 590850 444574 591430 444658
rect 590850 444338 591022 444574
rect 591258 444338 591430 444574
rect 590850 408894 591430 444338
rect 590850 408658 591022 408894
rect 591258 408658 591430 408894
rect 590850 408574 591430 408658
rect 590850 408338 591022 408574
rect 591258 408338 591430 408574
rect 590850 372894 591430 408338
rect 590850 372658 591022 372894
rect 591258 372658 591430 372894
rect 590850 372574 591430 372658
rect 590850 372338 591022 372574
rect 591258 372338 591430 372574
rect 590850 336894 591430 372338
rect 590850 336658 591022 336894
rect 591258 336658 591430 336894
rect 590850 336574 591430 336658
rect 590850 336338 591022 336574
rect 591258 336338 591430 336574
rect 590850 300894 591430 336338
rect 590850 300658 591022 300894
rect 591258 300658 591430 300894
rect 590850 300574 591430 300658
rect 590850 300338 591022 300574
rect 591258 300338 591430 300574
rect 590850 264894 591430 300338
rect 590850 264658 591022 264894
rect 591258 264658 591430 264894
rect 590850 264574 591430 264658
rect 590850 264338 591022 264574
rect 591258 264338 591430 264574
rect 590850 228894 591430 264338
rect 590850 228658 591022 228894
rect 591258 228658 591430 228894
rect 590850 228574 591430 228658
rect 590850 228338 591022 228574
rect 591258 228338 591430 228574
rect 590850 192894 591430 228338
rect 590850 192658 591022 192894
rect 591258 192658 591430 192894
rect 590850 192574 591430 192658
rect 590850 192338 591022 192574
rect 591258 192338 591430 192574
rect 590850 156894 591430 192338
rect 590850 156658 591022 156894
rect 591258 156658 591430 156894
rect 590850 156574 591430 156658
rect 590850 156338 591022 156574
rect 591258 156338 591430 156574
rect 590850 120894 591430 156338
rect 590850 120658 591022 120894
rect 591258 120658 591430 120894
rect 590850 120574 591430 120658
rect 590850 120338 591022 120574
rect 591258 120338 591430 120574
rect 590850 84894 591430 120338
rect 590850 84658 591022 84894
rect 591258 84658 591430 84894
rect 590850 84574 591430 84658
rect 590850 84338 591022 84574
rect 591258 84338 591430 84574
rect 590850 48894 591430 84338
rect 590850 48658 591022 48894
rect 591258 48658 591430 48894
rect 590850 48574 591430 48658
rect 590850 48338 591022 48574
rect 591258 48338 591430 48574
rect 590850 12894 591430 48338
rect 590850 12658 591022 12894
rect 591258 12658 591430 12894
rect 590850 12574 591430 12658
rect 590850 12338 591022 12574
rect 591258 12338 591430 12574
rect 590850 -5866 591430 12338
rect 590850 -6102 591022 -5866
rect 591258 -6102 591430 -5866
rect 590850 -6186 591430 -6102
rect 590850 -6422 591022 -6186
rect 591258 -6422 591430 -6186
rect 590850 -6434 591430 -6422
rect 591770 678894 592350 710722
rect 591770 678658 591942 678894
rect 592178 678658 592350 678894
rect 591770 678574 592350 678658
rect 591770 678338 591942 678574
rect 592178 678338 592350 678574
rect 591770 642894 592350 678338
rect 591770 642658 591942 642894
rect 592178 642658 592350 642894
rect 591770 642574 592350 642658
rect 591770 642338 591942 642574
rect 592178 642338 592350 642574
rect 591770 606894 592350 642338
rect 591770 606658 591942 606894
rect 592178 606658 592350 606894
rect 591770 606574 592350 606658
rect 591770 606338 591942 606574
rect 592178 606338 592350 606574
rect 591770 570894 592350 606338
rect 591770 570658 591942 570894
rect 592178 570658 592350 570894
rect 591770 570574 592350 570658
rect 591770 570338 591942 570574
rect 592178 570338 592350 570574
rect 591770 534894 592350 570338
rect 591770 534658 591942 534894
rect 592178 534658 592350 534894
rect 591770 534574 592350 534658
rect 591770 534338 591942 534574
rect 592178 534338 592350 534574
rect 591770 498894 592350 534338
rect 591770 498658 591942 498894
rect 592178 498658 592350 498894
rect 591770 498574 592350 498658
rect 591770 498338 591942 498574
rect 592178 498338 592350 498574
rect 591770 462894 592350 498338
rect 591770 462658 591942 462894
rect 592178 462658 592350 462894
rect 591770 462574 592350 462658
rect 591770 462338 591942 462574
rect 592178 462338 592350 462574
rect 591770 426894 592350 462338
rect 591770 426658 591942 426894
rect 592178 426658 592350 426894
rect 591770 426574 592350 426658
rect 591770 426338 591942 426574
rect 592178 426338 592350 426574
rect 591770 390894 592350 426338
rect 591770 390658 591942 390894
rect 592178 390658 592350 390894
rect 591770 390574 592350 390658
rect 591770 390338 591942 390574
rect 592178 390338 592350 390574
rect 591770 354894 592350 390338
rect 591770 354658 591942 354894
rect 592178 354658 592350 354894
rect 591770 354574 592350 354658
rect 591770 354338 591942 354574
rect 592178 354338 592350 354574
rect 591770 318894 592350 354338
rect 591770 318658 591942 318894
rect 592178 318658 592350 318894
rect 591770 318574 592350 318658
rect 591770 318338 591942 318574
rect 592178 318338 592350 318574
rect 591770 282894 592350 318338
rect 591770 282658 591942 282894
rect 592178 282658 592350 282894
rect 591770 282574 592350 282658
rect 591770 282338 591942 282574
rect 592178 282338 592350 282574
rect 591770 246894 592350 282338
rect 591770 246658 591942 246894
rect 592178 246658 592350 246894
rect 591770 246574 592350 246658
rect 591770 246338 591942 246574
rect 592178 246338 592350 246574
rect 591770 210894 592350 246338
rect 591770 210658 591942 210894
rect 592178 210658 592350 210894
rect 591770 210574 592350 210658
rect 591770 210338 591942 210574
rect 592178 210338 592350 210574
rect 591770 174894 592350 210338
rect 591770 174658 591942 174894
rect 592178 174658 592350 174894
rect 591770 174574 592350 174658
rect 591770 174338 591942 174574
rect 592178 174338 592350 174574
rect 591770 138894 592350 174338
rect 591770 138658 591942 138894
rect 592178 138658 592350 138894
rect 591770 138574 592350 138658
rect 591770 138338 591942 138574
rect 592178 138338 592350 138574
rect 591770 102894 592350 138338
rect 591770 102658 591942 102894
rect 592178 102658 592350 102894
rect 591770 102574 592350 102658
rect 591770 102338 591942 102574
rect 592178 102338 592350 102574
rect 591770 66894 592350 102338
rect 591770 66658 591942 66894
rect 592178 66658 592350 66894
rect 591770 66574 592350 66658
rect 591770 66338 591942 66574
rect 592178 66338 592350 66574
rect 591770 30894 592350 66338
rect 591770 30658 591942 30894
rect 592178 30658 592350 30894
rect 591770 30574 592350 30658
rect 591770 30338 591942 30574
rect 592178 30338 592350 30574
rect 569254 -7022 569426 -6786
rect 569662 -7022 569834 -6786
rect 569254 -7106 569834 -7022
rect 569254 -7342 569426 -7106
rect 569662 -7342 569834 -7106
rect 569254 -7354 569834 -7342
rect 591770 -6786 592350 30338
rect 591770 -7022 591942 -6786
rect 592178 -7022 592350 -6786
rect 591770 -7106 592350 -7022
rect 591770 -7342 591942 -7106
rect 592178 -7342 592350 -7106
rect 591770 -7354 592350 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 678658 -8018 678894
rect -8254 678338 -8018 678574
rect -8254 642658 -8018 642894
rect -8254 642338 -8018 642574
rect -8254 606658 -8018 606894
rect -8254 606338 -8018 606574
rect -8254 570658 -8018 570894
rect -8254 570338 -8018 570574
rect -8254 534658 -8018 534894
rect -8254 534338 -8018 534574
rect -8254 498658 -8018 498894
rect -8254 498338 -8018 498574
rect -8254 462658 -8018 462894
rect -8254 462338 -8018 462574
rect -8254 426658 -8018 426894
rect -8254 426338 -8018 426574
rect -8254 390658 -8018 390894
rect -8254 390338 -8018 390574
rect -8254 354658 -8018 354894
rect -8254 354338 -8018 354574
rect -8254 318658 -8018 318894
rect -8254 318338 -8018 318574
rect -8254 282658 -8018 282894
rect -8254 282338 -8018 282574
rect -8254 246658 -8018 246894
rect -8254 246338 -8018 246574
rect -8254 210658 -8018 210894
rect -8254 210338 -8018 210574
rect -8254 174658 -8018 174894
rect -8254 174338 -8018 174574
rect -8254 138658 -8018 138894
rect -8254 138338 -8018 138574
rect -8254 102658 -8018 102894
rect -8254 102338 -8018 102574
rect -8254 66658 -8018 66894
rect -8254 66338 -8018 66574
rect -8254 30658 -8018 30894
rect -8254 30338 -8018 30574
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11426 710122 11662 710358
rect 11426 709802 11662 710038
rect -7334 696658 -7098 696894
rect -7334 696338 -7098 696574
rect -7334 660658 -7098 660894
rect -7334 660338 -7098 660574
rect -7334 624658 -7098 624894
rect -7334 624338 -7098 624574
rect -7334 588658 -7098 588894
rect -7334 588338 -7098 588574
rect -7334 552658 -7098 552894
rect -7334 552338 -7098 552574
rect -7334 516658 -7098 516894
rect -7334 516338 -7098 516574
rect -7334 480658 -7098 480894
rect -7334 480338 -7098 480574
rect -7334 444658 -7098 444894
rect -7334 444338 -7098 444574
rect -7334 408658 -7098 408894
rect -7334 408338 -7098 408574
rect -7334 372658 -7098 372894
rect -7334 372338 -7098 372574
rect -7334 336658 -7098 336894
rect -7334 336338 -7098 336574
rect -7334 300658 -7098 300894
rect -7334 300338 -7098 300574
rect -7334 264658 -7098 264894
rect -7334 264338 -7098 264574
rect -7334 228658 -7098 228894
rect -7334 228338 -7098 228574
rect -7334 192658 -7098 192894
rect -7334 192338 -7098 192574
rect -7334 156658 -7098 156894
rect -7334 156338 -7098 156574
rect -7334 120658 -7098 120894
rect -7334 120338 -7098 120574
rect -7334 84658 -7098 84894
rect -7334 84338 -7098 84574
rect -7334 48658 -7098 48894
rect -7334 48338 -7098 48574
rect -7334 12658 -7098 12894
rect -7334 12338 -7098 12574
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675178 -6178 675414
rect -6414 674858 -6178 675094
rect -6414 639178 -6178 639414
rect -6414 638858 -6178 639094
rect -6414 603178 -6178 603414
rect -6414 602858 -6178 603094
rect -6414 567178 -6178 567414
rect -6414 566858 -6178 567094
rect -6414 531178 -6178 531414
rect -6414 530858 -6178 531094
rect -6414 495178 -6178 495414
rect -6414 494858 -6178 495094
rect -6414 459178 -6178 459414
rect -6414 458858 -6178 459094
rect -6414 423178 -6178 423414
rect -6414 422858 -6178 423094
rect -6414 387178 -6178 387414
rect -6414 386858 -6178 387094
rect -6414 351178 -6178 351414
rect -6414 350858 -6178 351094
rect -6414 315178 -6178 315414
rect -6414 314858 -6178 315094
rect -6414 279178 -6178 279414
rect -6414 278858 -6178 279094
rect -6414 243178 -6178 243414
rect -6414 242858 -6178 243094
rect -6414 207178 -6178 207414
rect -6414 206858 -6178 207094
rect -6414 171178 -6178 171414
rect -6414 170858 -6178 171094
rect -6414 135178 -6178 135414
rect -6414 134858 -6178 135094
rect -6414 99178 -6178 99414
rect -6414 98858 -6178 99094
rect -6414 63178 -6178 63414
rect -6414 62858 -6178 63094
rect -6414 27178 -6178 27414
rect -6414 26858 -6178 27094
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 7946 708282 8182 708518
rect 7946 707962 8182 708198
rect -5494 693178 -5258 693414
rect -5494 692858 -5258 693094
rect -5494 657178 -5258 657414
rect -5494 656858 -5258 657094
rect -5494 621178 -5258 621414
rect -5494 620858 -5258 621094
rect -5494 585178 -5258 585414
rect -5494 584858 -5258 585094
rect -5494 549178 -5258 549414
rect -5494 548858 -5258 549094
rect -5494 513178 -5258 513414
rect -5494 512858 -5258 513094
rect -5494 477178 -5258 477414
rect -5494 476858 -5258 477094
rect -5494 441178 -5258 441414
rect -5494 440858 -5258 441094
rect -5494 405178 -5258 405414
rect -5494 404858 -5258 405094
rect -5494 369178 -5258 369414
rect -5494 368858 -5258 369094
rect -5494 333178 -5258 333414
rect -5494 332858 -5258 333094
rect -5494 297178 -5258 297414
rect -5494 296858 -5258 297094
rect -5494 261178 -5258 261414
rect -5494 260858 -5258 261094
rect -5494 225178 -5258 225414
rect -5494 224858 -5258 225094
rect -5494 189178 -5258 189414
rect -5494 188858 -5258 189094
rect -5494 153178 -5258 153414
rect -5494 152858 -5258 153094
rect -5494 117178 -5258 117414
rect -5494 116858 -5258 117094
rect -5494 81178 -5258 81414
rect -5494 80858 -5258 81094
rect -5494 45178 -5258 45414
rect -5494 44858 -5258 45094
rect -5494 9178 -5258 9414
rect -5494 8858 -5258 9094
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671698 -4338 671934
rect -4574 671378 -4338 671614
rect -4574 635698 -4338 635934
rect -4574 635378 -4338 635614
rect -4574 599698 -4338 599934
rect -4574 599378 -4338 599614
rect -4574 563698 -4338 563934
rect -4574 563378 -4338 563614
rect -4574 527698 -4338 527934
rect -4574 527378 -4338 527614
rect -4574 491698 -4338 491934
rect -4574 491378 -4338 491614
rect -4574 455698 -4338 455934
rect -4574 455378 -4338 455614
rect -4574 419698 -4338 419934
rect -4574 419378 -4338 419614
rect -4574 383698 -4338 383934
rect -4574 383378 -4338 383614
rect -4574 347698 -4338 347934
rect -4574 347378 -4338 347614
rect -4574 311698 -4338 311934
rect -4574 311378 -4338 311614
rect -4574 275698 -4338 275934
rect -4574 275378 -4338 275614
rect -4574 239698 -4338 239934
rect -4574 239378 -4338 239614
rect -4574 203698 -4338 203934
rect -4574 203378 -4338 203614
rect -4574 167698 -4338 167934
rect -4574 167378 -4338 167614
rect -4574 131698 -4338 131934
rect -4574 131378 -4338 131614
rect -4574 95698 -4338 95934
rect -4574 95378 -4338 95614
rect -4574 59698 -4338 59934
rect -4574 59378 -4338 59614
rect -4574 23698 -4338 23934
rect -4574 23378 -4338 23614
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4466 706442 4702 706678
rect 4466 706122 4702 706358
rect -3654 689698 -3418 689934
rect -3654 689378 -3418 689614
rect -3654 653698 -3418 653934
rect -3654 653378 -3418 653614
rect -3654 617698 -3418 617934
rect -3654 617378 -3418 617614
rect -3654 581698 -3418 581934
rect -3654 581378 -3418 581614
rect -3654 545698 -3418 545934
rect -3654 545378 -3418 545614
rect -3654 509698 -3418 509934
rect -3654 509378 -3418 509614
rect -3654 473698 -3418 473934
rect -3654 473378 -3418 473614
rect -3654 437698 -3418 437934
rect -3654 437378 -3418 437614
rect -3654 401698 -3418 401934
rect -3654 401378 -3418 401614
rect -3654 365698 -3418 365934
rect -3654 365378 -3418 365614
rect -3654 329698 -3418 329934
rect -3654 329378 -3418 329614
rect -3654 293698 -3418 293934
rect -3654 293378 -3418 293614
rect -3654 257698 -3418 257934
rect -3654 257378 -3418 257614
rect -3654 221698 -3418 221934
rect -3654 221378 -3418 221614
rect -3654 185698 -3418 185934
rect -3654 185378 -3418 185614
rect -3654 149698 -3418 149934
rect -3654 149378 -3418 149614
rect -3654 113698 -3418 113934
rect -3654 113378 -3418 113614
rect -3654 77698 -3418 77934
rect -3654 77378 -3418 77614
rect -3654 41698 -3418 41934
rect -3654 41378 -3418 41614
rect -3654 5698 -3418 5934
rect -3654 5378 -3418 5614
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4466 689698 4702 689934
rect 4466 689378 4702 689614
rect 4466 653698 4702 653934
rect 4466 653378 4702 653614
rect 4466 617698 4702 617934
rect 4466 617378 4702 617614
rect 4466 581698 4702 581934
rect 4466 581378 4702 581614
rect 4466 545698 4702 545934
rect 4466 545378 4702 545614
rect 4466 509698 4702 509934
rect 4466 509378 4702 509614
rect 4466 473698 4702 473934
rect 4466 473378 4702 473614
rect 4466 437698 4702 437934
rect 4466 437378 4702 437614
rect 4466 401698 4702 401934
rect 4466 401378 4702 401614
rect 4466 365698 4702 365934
rect 4466 365378 4702 365614
rect 4466 329698 4702 329934
rect 4466 329378 4702 329614
rect 4466 293698 4702 293934
rect 4466 293378 4702 293614
rect 4466 257698 4702 257934
rect 4466 257378 4702 257614
rect 4466 221698 4702 221934
rect 4466 221378 4702 221614
rect 4466 185698 4702 185934
rect 4466 185378 4702 185614
rect 4466 149698 4702 149934
rect 4466 149378 4702 149614
rect 4466 113698 4702 113934
rect 4466 113378 4702 113614
rect 4466 77698 4702 77934
rect 4466 77378 4702 77614
rect 4466 41698 4702 41934
rect 4466 41378 4702 41614
rect 4466 5698 4702 5934
rect 4466 5378 4702 5614
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4466 -2422 4702 -2186
rect 4466 -2742 4702 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 7946 693178 8182 693414
rect 7946 692858 8182 693094
rect 7946 657178 8182 657414
rect 7946 656858 8182 657094
rect 7946 621178 8182 621414
rect 7946 620858 8182 621094
rect 7946 585178 8182 585414
rect 7946 584858 8182 585094
rect 7946 549178 8182 549414
rect 7946 548858 8182 549094
rect 7946 513178 8182 513414
rect 7946 512858 8182 513094
rect 7946 477178 8182 477414
rect 7946 476858 8182 477094
rect 7946 441178 8182 441414
rect 7946 440858 8182 441094
rect 7946 405178 8182 405414
rect 7946 404858 8182 405094
rect 7946 369178 8182 369414
rect 7946 368858 8182 369094
rect 7946 333178 8182 333414
rect 7946 332858 8182 333094
rect 7946 297178 8182 297414
rect 7946 296858 8182 297094
rect 7946 261178 8182 261414
rect 7946 260858 8182 261094
rect 7946 225178 8182 225414
rect 7946 224858 8182 225094
rect 7946 189178 8182 189414
rect 7946 188858 8182 189094
rect 7946 153178 8182 153414
rect 7946 152858 8182 153094
rect 7946 117178 8182 117414
rect 7946 116858 8182 117094
rect 7946 81178 8182 81414
rect 7946 80858 8182 81094
rect 7946 45178 8182 45414
rect 7946 44858 8182 45094
rect 7946 9178 8182 9414
rect 7946 8858 8182 9094
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 7946 -4262 8182 -4026
rect 7946 -4582 8182 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29426 711042 29662 711278
rect 29426 710722 29662 710958
rect 25946 709202 26182 709438
rect 25946 708882 26182 709118
rect 22466 707362 22702 707598
rect 22466 707042 22702 707278
rect 11426 696658 11662 696894
rect 11426 696338 11662 696574
rect 11426 660658 11662 660894
rect 11426 660338 11662 660574
rect 11426 624658 11662 624894
rect 11426 624338 11662 624574
rect 11426 588658 11662 588894
rect 11426 588338 11662 588574
rect 11426 552658 11662 552894
rect 11426 552338 11662 552574
rect 11426 516658 11662 516894
rect 11426 516338 11662 516574
rect 11426 480658 11662 480894
rect 11426 480338 11662 480574
rect 11426 444658 11662 444894
rect 11426 444338 11662 444574
rect 11426 408658 11662 408894
rect 11426 408338 11662 408574
rect 11426 372658 11662 372894
rect 11426 372338 11662 372574
rect 11426 336658 11662 336894
rect 11426 336338 11662 336574
rect 11426 300658 11662 300894
rect 11426 300338 11662 300574
rect 11426 264658 11662 264894
rect 11426 264338 11662 264574
rect 11426 228658 11662 228894
rect 11426 228338 11662 228574
rect 11426 192658 11662 192894
rect 11426 192338 11662 192574
rect 11426 156658 11662 156894
rect 11426 156338 11662 156574
rect 11426 120658 11662 120894
rect 11426 120338 11662 120574
rect 11426 84658 11662 84894
rect 11426 84338 11662 84574
rect 11426 48658 11662 48894
rect 11426 48338 11662 48574
rect 11426 12658 11662 12894
rect 11426 12338 11662 12574
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22466 671698 22702 671934
rect 22466 671378 22702 671614
rect 22466 635698 22702 635934
rect 22466 635378 22702 635614
rect 22466 599698 22702 599934
rect 22466 599378 22702 599614
rect 22466 563698 22702 563934
rect 22466 563378 22702 563614
rect 22466 527698 22702 527934
rect 22466 527378 22702 527614
rect 22466 491698 22702 491934
rect 22466 491378 22702 491614
rect 22466 455698 22702 455934
rect 22466 455378 22702 455614
rect 22466 419698 22702 419934
rect 22466 419378 22702 419614
rect 22466 383698 22702 383934
rect 22466 383378 22702 383614
rect 22466 347698 22702 347934
rect 22466 347378 22702 347614
rect 22466 311698 22702 311934
rect 22466 311378 22702 311614
rect 22466 275698 22702 275934
rect 22466 275378 22702 275614
rect 22466 239698 22702 239934
rect 22466 239378 22702 239614
rect 22466 203698 22702 203934
rect 22466 203378 22702 203614
rect 22466 167698 22702 167934
rect 22466 167378 22702 167614
rect 22466 131698 22702 131934
rect 22466 131378 22702 131614
rect 22466 95698 22702 95934
rect 22466 95378 22702 95614
rect 22466 59698 22702 59934
rect 22466 59378 22702 59614
rect 22466 23698 22702 23934
rect 22466 23378 22702 23614
rect 22466 -3342 22702 -3106
rect 22466 -3662 22702 -3426
rect 25946 675178 26182 675414
rect 25946 674858 26182 675094
rect 25946 639178 26182 639414
rect 25946 638858 26182 639094
rect 25946 603178 26182 603414
rect 25946 602858 26182 603094
rect 25946 567178 26182 567414
rect 25946 566858 26182 567094
rect 25946 531178 26182 531414
rect 25946 530858 26182 531094
rect 25946 495178 26182 495414
rect 25946 494858 26182 495094
rect 25946 459178 26182 459414
rect 25946 458858 26182 459094
rect 25946 423178 26182 423414
rect 25946 422858 26182 423094
rect 25946 387178 26182 387414
rect 25946 386858 26182 387094
rect 25946 351178 26182 351414
rect 25946 350858 26182 351094
rect 25946 315178 26182 315414
rect 25946 314858 26182 315094
rect 25946 279178 26182 279414
rect 25946 278858 26182 279094
rect 25946 243178 26182 243414
rect 25946 242858 26182 243094
rect 25946 207178 26182 207414
rect 25946 206858 26182 207094
rect 25946 171178 26182 171414
rect 25946 170858 26182 171094
rect 25946 135178 26182 135414
rect 25946 134858 26182 135094
rect 25946 99178 26182 99414
rect 25946 98858 26182 99094
rect 25946 63178 26182 63414
rect 25946 62858 26182 63094
rect 25946 27178 26182 27414
rect 25946 26858 26182 27094
rect 25946 -5182 26182 -4946
rect 25946 -5502 26182 -5266
rect 47426 710122 47662 710358
rect 47426 709802 47662 710038
rect 43946 708282 44182 708518
rect 43946 707962 44182 708198
rect 40466 706442 40702 706678
rect 40466 706122 40702 706358
rect 29426 678658 29662 678894
rect 29426 678338 29662 678574
rect 29426 642658 29662 642894
rect 29426 642338 29662 642574
rect 29426 606658 29662 606894
rect 29426 606338 29662 606574
rect 29426 570658 29662 570894
rect 29426 570338 29662 570574
rect 29426 534658 29662 534894
rect 29426 534338 29662 534574
rect 29426 498658 29662 498894
rect 29426 498338 29662 498574
rect 29426 462658 29662 462894
rect 29426 462338 29662 462574
rect 29426 426658 29662 426894
rect 29426 426338 29662 426574
rect 29426 390658 29662 390894
rect 29426 390338 29662 390574
rect 29426 354658 29662 354894
rect 29426 354338 29662 354574
rect 29426 318658 29662 318894
rect 29426 318338 29662 318574
rect 29426 282658 29662 282894
rect 29426 282338 29662 282574
rect 29426 246658 29662 246894
rect 29426 246338 29662 246574
rect 29426 210658 29662 210894
rect 29426 210338 29662 210574
rect 29426 174658 29662 174894
rect 29426 174338 29662 174574
rect 29426 138658 29662 138894
rect 29426 138338 29662 138574
rect 29426 102658 29662 102894
rect 29426 102338 29662 102574
rect 29426 66658 29662 66894
rect 29426 66338 29662 66574
rect 29426 30658 29662 30894
rect 29426 30338 29662 30574
rect 11426 -6102 11662 -5866
rect 11426 -6422 11662 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40466 689698 40702 689934
rect 40466 689378 40702 689614
rect 40466 653698 40702 653934
rect 40466 653378 40702 653614
rect 40466 617698 40702 617934
rect 40466 617378 40702 617614
rect 40466 581698 40702 581934
rect 40466 581378 40702 581614
rect 40466 545698 40702 545934
rect 40466 545378 40702 545614
rect 40466 509698 40702 509934
rect 40466 509378 40702 509614
rect 40466 473698 40702 473934
rect 40466 473378 40702 473614
rect 40466 437698 40702 437934
rect 40466 437378 40702 437614
rect 40466 401698 40702 401934
rect 40466 401378 40702 401614
rect 40466 365698 40702 365934
rect 40466 365378 40702 365614
rect 40466 329698 40702 329934
rect 40466 329378 40702 329614
rect 40466 293698 40702 293934
rect 40466 293378 40702 293614
rect 40466 257698 40702 257934
rect 40466 257378 40702 257614
rect 40466 221698 40702 221934
rect 40466 221378 40702 221614
rect 40466 185698 40702 185934
rect 40466 185378 40702 185614
rect 40466 149698 40702 149934
rect 40466 149378 40702 149614
rect 40466 113698 40702 113934
rect 40466 113378 40702 113614
rect 40466 77698 40702 77934
rect 40466 77378 40702 77614
rect 40466 41698 40702 41934
rect 40466 41378 40702 41614
rect 40466 5698 40702 5934
rect 40466 5378 40702 5614
rect 40466 -2422 40702 -2186
rect 40466 -2742 40702 -2506
rect 43946 693178 44182 693414
rect 43946 692858 44182 693094
rect 43946 657178 44182 657414
rect 43946 656858 44182 657094
rect 43946 621178 44182 621414
rect 43946 620858 44182 621094
rect 43946 585178 44182 585414
rect 43946 584858 44182 585094
rect 43946 549178 44182 549414
rect 43946 548858 44182 549094
rect 43946 513178 44182 513414
rect 43946 512858 44182 513094
rect 43946 477178 44182 477414
rect 43946 476858 44182 477094
rect 43946 441178 44182 441414
rect 43946 440858 44182 441094
rect 43946 405178 44182 405414
rect 43946 404858 44182 405094
rect 43946 369178 44182 369414
rect 43946 368858 44182 369094
rect 43946 333178 44182 333414
rect 43946 332858 44182 333094
rect 43946 297178 44182 297414
rect 43946 296858 44182 297094
rect 43946 261178 44182 261414
rect 43946 260858 44182 261094
rect 43946 225178 44182 225414
rect 43946 224858 44182 225094
rect 43946 189178 44182 189414
rect 43946 188858 44182 189094
rect 43946 153178 44182 153414
rect 43946 152858 44182 153094
rect 43946 117178 44182 117414
rect 43946 116858 44182 117094
rect 43946 81178 44182 81414
rect 43946 80858 44182 81094
rect 43946 45178 44182 45414
rect 43946 44858 44182 45094
rect 43946 9178 44182 9414
rect 43946 8858 44182 9094
rect 43946 -4262 44182 -4026
rect 43946 -4582 44182 -4346
rect 65426 711042 65662 711278
rect 65426 710722 65662 710958
rect 61946 709202 62182 709438
rect 61946 708882 62182 709118
rect 58466 707362 58702 707598
rect 58466 707042 58702 707278
rect 47426 696658 47662 696894
rect 47426 696338 47662 696574
rect 47426 660658 47662 660894
rect 47426 660338 47662 660574
rect 47426 624658 47662 624894
rect 47426 624338 47662 624574
rect 47426 588658 47662 588894
rect 47426 588338 47662 588574
rect 47426 552658 47662 552894
rect 47426 552338 47662 552574
rect 47426 516658 47662 516894
rect 47426 516338 47662 516574
rect 47426 480658 47662 480894
rect 47426 480338 47662 480574
rect 47426 444658 47662 444894
rect 47426 444338 47662 444574
rect 47426 408658 47662 408894
rect 47426 408338 47662 408574
rect 47426 372658 47662 372894
rect 47426 372338 47662 372574
rect 47426 336658 47662 336894
rect 47426 336338 47662 336574
rect 47426 300658 47662 300894
rect 47426 300338 47662 300574
rect 47426 264658 47662 264894
rect 47426 264338 47662 264574
rect 47426 228658 47662 228894
rect 47426 228338 47662 228574
rect 47426 192658 47662 192894
rect 47426 192338 47662 192574
rect 47426 156658 47662 156894
rect 47426 156338 47662 156574
rect 47426 120658 47662 120894
rect 47426 120338 47662 120574
rect 47426 84658 47662 84894
rect 47426 84338 47662 84574
rect 47426 48658 47662 48894
rect 47426 48338 47662 48574
rect 47426 12658 47662 12894
rect 47426 12338 47662 12574
rect 29426 -7022 29662 -6786
rect 29426 -7342 29662 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58466 671698 58702 671934
rect 58466 671378 58702 671614
rect 58466 635698 58702 635934
rect 58466 635378 58702 635614
rect 58466 599698 58702 599934
rect 58466 599378 58702 599614
rect 58466 563698 58702 563934
rect 58466 563378 58702 563614
rect 58466 527698 58702 527934
rect 58466 527378 58702 527614
rect 58466 491698 58702 491934
rect 58466 491378 58702 491614
rect 58466 455698 58702 455934
rect 58466 455378 58702 455614
rect 58466 419698 58702 419934
rect 58466 419378 58702 419614
rect 58466 383698 58702 383934
rect 58466 383378 58702 383614
rect 58466 347698 58702 347934
rect 58466 347378 58702 347614
rect 58466 311698 58702 311934
rect 58466 311378 58702 311614
rect 58466 275698 58702 275934
rect 58466 275378 58702 275614
rect 58466 239698 58702 239934
rect 58466 239378 58702 239614
rect 58466 203698 58702 203934
rect 58466 203378 58702 203614
rect 58466 167698 58702 167934
rect 58466 167378 58702 167614
rect 58466 131698 58702 131934
rect 58466 131378 58702 131614
rect 58466 95698 58702 95934
rect 58466 95378 58702 95614
rect 58466 59698 58702 59934
rect 58466 59378 58702 59614
rect 58466 23698 58702 23934
rect 58466 23378 58702 23614
rect 58466 -3342 58702 -3106
rect 58466 -3662 58702 -3426
rect 61946 675178 62182 675414
rect 61946 674858 62182 675094
rect 61946 639178 62182 639414
rect 61946 638858 62182 639094
rect 61946 603178 62182 603414
rect 61946 602858 62182 603094
rect 61946 567178 62182 567414
rect 61946 566858 62182 567094
rect 61946 531178 62182 531414
rect 61946 530858 62182 531094
rect 61946 495178 62182 495414
rect 61946 494858 62182 495094
rect 61946 459178 62182 459414
rect 61946 458858 62182 459094
rect 61946 423178 62182 423414
rect 61946 422858 62182 423094
rect 61946 387178 62182 387414
rect 61946 386858 62182 387094
rect 61946 351178 62182 351414
rect 61946 350858 62182 351094
rect 61946 315178 62182 315414
rect 61946 314858 62182 315094
rect 61946 279178 62182 279414
rect 61946 278858 62182 279094
rect 61946 243178 62182 243414
rect 61946 242858 62182 243094
rect 61946 207178 62182 207414
rect 61946 206858 62182 207094
rect 61946 171178 62182 171414
rect 61946 170858 62182 171094
rect 61946 135178 62182 135414
rect 61946 134858 62182 135094
rect 61946 99178 62182 99414
rect 61946 98858 62182 99094
rect 61946 63178 62182 63414
rect 61946 62858 62182 63094
rect 61946 27178 62182 27414
rect 61946 26858 62182 27094
rect 61946 -5182 62182 -4946
rect 61946 -5502 62182 -5266
rect 83426 710122 83662 710358
rect 83426 709802 83662 710038
rect 79946 708282 80182 708518
rect 79946 707962 80182 708198
rect 76466 706442 76702 706678
rect 76466 706122 76702 706358
rect 65426 678658 65662 678894
rect 65426 678338 65662 678574
rect 65426 642658 65662 642894
rect 65426 642338 65662 642574
rect 65426 606658 65662 606894
rect 65426 606338 65662 606574
rect 65426 570658 65662 570894
rect 65426 570338 65662 570574
rect 65426 534658 65662 534894
rect 65426 534338 65662 534574
rect 65426 498658 65662 498894
rect 65426 498338 65662 498574
rect 65426 462658 65662 462894
rect 65426 462338 65662 462574
rect 65426 426658 65662 426894
rect 65426 426338 65662 426574
rect 65426 390658 65662 390894
rect 65426 390338 65662 390574
rect 65426 354658 65662 354894
rect 65426 354338 65662 354574
rect 65426 318658 65662 318894
rect 65426 318338 65662 318574
rect 65426 282658 65662 282894
rect 65426 282338 65662 282574
rect 65426 246658 65662 246894
rect 65426 246338 65662 246574
rect 65426 210658 65662 210894
rect 65426 210338 65662 210574
rect 65426 174658 65662 174894
rect 65426 174338 65662 174574
rect 65426 138658 65662 138894
rect 65426 138338 65662 138574
rect 65426 102658 65662 102894
rect 65426 102338 65662 102574
rect 65426 66658 65662 66894
rect 65426 66338 65662 66574
rect 65426 30658 65662 30894
rect 65426 30338 65662 30574
rect 47426 -6102 47662 -5866
rect 47426 -6422 47662 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76466 689698 76702 689934
rect 76466 689378 76702 689614
rect 76466 653698 76702 653934
rect 76466 653378 76702 653614
rect 76466 617698 76702 617934
rect 76466 617378 76702 617614
rect 76466 581698 76702 581934
rect 76466 581378 76702 581614
rect 76466 545698 76702 545934
rect 76466 545378 76702 545614
rect 76466 509698 76702 509934
rect 76466 509378 76702 509614
rect 76466 473698 76702 473934
rect 76466 473378 76702 473614
rect 76466 437698 76702 437934
rect 76466 437378 76702 437614
rect 76466 401698 76702 401934
rect 76466 401378 76702 401614
rect 76466 365698 76702 365934
rect 76466 365378 76702 365614
rect 76466 329698 76702 329934
rect 76466 329378 76702 329614
rect 76466 293698 76702 293934
rect 76466 293378 76702 293614
rect 76466 257698 76702 257934
rect 76466 257378 76702 257614
rect 76466 221698 76702 221934
rect 76466 221378 76702 221614
rect 76466 185698 76702 185934
rect 76466 185378 76702 185614
rect 76466 149698 76702 149934
rect 76466 149378 76702 149614
rect 76466 113698 76702 113934
rect 76466 113378 76702 113614
rect 76466 77698 76702 77934
rect 76466 77378 76702 77614
rect 76466 41698 76702 41934
rect 76466 41378 76702 41614
rect 76466 5698 76702 5934
rect 76466 5378 76702 5614
rect 76466 -2422 76702 -2186
rect 76466 -2742 76702 -2506
rect 79946 693178 80182 693414
rect 79946 692858 80182 693094
rect 79946 657178 80182 657414
rect 79946 656858 80182 657094
rect 79946 621178 80182 621414
rect 79946 620858 80182 621094
rect 79946 585178 80182 585414
rect 79946 584858 80182 585094
rect 79946 549178 80182 549414
rect 79946 548858 80182 549094
rect 79946 513178 80182 513414
rect 79946 512858 80182 513094
rect 79946 477178 80182 477414
rect 79946 476858 80182 477094
rect 79946 441178 80182 441414
rect 79946 440858 80182 441094
rect 79946 405178 80182 405414
rect 79946 404858 80182 405094
rect 79946 369178 80182 369414
rect 79946 368858 80182 369094
rect 79946 333178 80182 333414
rect 79946 332858 80182 333094
rect 79946 297178 80182 297414
rect 79946 296858 80182 297094
rect 79946 261178 80182 261414
rect 79946 260858 80182 261094
rect 79946 225178 80182 225414
rect 79946 224858 80182 225094
rect 79946 189178 80182 189414
rect 79946 188858 80182 189094
rect 79946 153178 80182 153414
rect 79946 152858 80182 153094
rect 79946 117178 80182 117414
rect 79946 116858 80182 117094
rect 79946 81178 80182 81414
rect 79946 80858 80182 81094
rect 79946 45178 80182 45414
rect 79946 44858 80182 45094
rect 79946 9178 80182 9414
rect 79946 8858 80182 9094
rect 79946 -4262 80182 -4026
rect 79946 -4582 80182 -4346
rect 101426 711042 101662 711278
rect 101426 710722 101662 710958
rect 97946 709202 98182 709438
rect 97946 708882 98182 709118
rect 94466 707362 94702 707598
rect 94466 707042 94702 707278
rect 83426 696658 83662 696894
rect 83426 696338 83662 696574
rect 83426 660658 83662 660894
rect 83426 660338 83662 660574
rect 83426 624658 83662 624894
rect 83426 624338 83662 624574
rect 83426 588658 83662 588894
rect 83426 588338 83662 588574
rect 83426 552658 83662 552894
rect 83426 552338 83662 552574
rect 83426 516658 83662 516894
rect 83426 516338 83662 516574
rect 83426 480658 83662 480894
rect 83426 480338 83662 480574
rect 83426 444658 83662 444894
rect 83426 444338 83662 444574
rect 83426 408658 83662 408894
rect 83426 408338 83662 408574
rect 83426 372658 83662 372894
rect 83426 372338 83662 372574
rect 83426 336658 83662 336894
rect 83426 336338 83662 336574
rect 83426 300658 83662 300894
rect 83426 300338 83662 300574
rect 83426 264658 83662 264894
rect 83426 264338 83662 264574
rect 83426 228658 83662 228894
rect 83426 228338 83662 228574
rect 83426 192658 83662 192894
rect 83426 192338 83662 192574
rect 83426 156658 83662 156894
rect 83426 156338 83662 156574
rect 83426 120658 83662 120894
rect 83426 120338 83662 120574
rect 83426 84658 83662 84894
rect 83426 84338 83662 84574
rect 83426 48658 83662 48894
rect 83426 48338 83662 48574
rect 83426 12658 83662 12894
rect 83426 12338 83662 12574
rect 65426 -7022 65662 -6786
rect 65426 -7342 65662 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94466 671698 94702 671934
rect 94466 671378 94702 671614
rect 94466 635698 94702 635934
rect 94466 635378 94702 635614
rect 94466 599698 94702 599934
rect 94466 599378 94702 599614
rect 94466 563698 94702 563934
rect 94466 563378 94702 563614
rect 94466 527698 94702 527934
rect 94466 527378 94702 527614
rect 94466 491698 94702 491934
rect 94466 491378 94702 491614
rect 94466 455698 94702 455934
rect 94466 455378 94702 455614
rect 94466 419698 94702 419934
rect 94466 419378 94702 419614
rect 94466 383698 94702 383934
rect 94466 383378 94702 383614
rect 94466 347698 94702 347934
rect 94466 347378 94702 347614
rect 94466 311698 94702 311934
rect 94466 311378 94702 311614
rect 94466 275698 94702 275934
rect 94466 275378 94702 275614
rect 94466 239698 94702 239934
rect 94466 239378 94702 239614
rect 94466 203698 94702 203934
rect 94466 203378 94702 203614
rect 94466 167698 94702 167934
rect 94466 167378 94702 167614
rect 94466 131698 94702 131934
rect 94466 131378 94702 131614
rect 94466 95698 94702 95934
rect 94466 95378 94702 95614
rect 94466 59698 94702 59934
rect 94466 59378 94702 59614
rect 94466 23698 94702 23934
rect 94466 23378 94702 23614
rect 94466 -3342 94702 -3106
rect 94466 -3662 94702 -3426
rect 97946 675178 98182 675414
rect 97946 674858 98182 675094
rect 97946 639178 98182 639414
rect 97946 638858 98182 639094
rect 97946 603178 98182 603414
rect 97946 602858 98182 603094
rect 97946 567178 98182 567414
rect 97946 566858 98182 567094
rect 97946 531178 98182 531414
rect 97946 530858 98182 531094
rect 97946 495178 98182 495414
rect 97946 494858 98182 495094
rect 97946 459178 98182 459414
rect 97946 458858 98182 459094
rect 97946 423178 98182 423414
rect 97946 422858 98182 423094
rect 97946 387178 98182 387414
rect 97946 386858 98182 387094
rect 97946 351178 98182 351414
rect 97946 350858 98182 351094
rect 97946 315178 98182 315414
rect 97946 314858 98182 315094
rect 97946 279178 98182 279414
rect 97946 278858 98182 279094
rect 97946 243178 98182 243414
rect 97946 242858 98182 243094
rect 97946 207178 98182 207414
rect 97946 206858 98182 207094
rect 97946 171178 98182 171414
rect 97946 170858 98182 171094
rect 97946 135178 98182 135414
rect 97946 134858 98182 135094
rect 97946 99178 98182 99414
rect 97946 98858 98182 99094
rect 97946 63178 98182 63414
rect 97946 62858 98182 63094
rect 97946 27178 98182 27414
rect 97946 26858 98182 27094
rect 97946 -5182 98182 -4946
rect 97946 -5502 98182 -5266
rect 119426 710122 119662 710358
rect 119426 709802 119662 710038
rect 115946 708282 116182 708518
rect 115946 707962 116182 708198
rect 112466 706442 112702 706678
rect 112466 706122 112702 706358
rect 101426 678658 101662 678894
rect 101426 678338 101662 678574
rect 101426 642658 101662 642894
rect 101426 642338 101662 642574
rect 101426 606658 101662 606894
rect 101426 606338 101662 606574
rect 101426 570658 101662 570894
rect 101426 570338 101662 570574
rect 101426 534658 101662 534894
rect 101426 534338 101662 534574
rect 101426 498658 101662 498894
rect 101426 498338 101662 498574
rect 101426 462658 101662 462894
rect 101426 462338 101662 462574
rect 101426 426658 101662 426894
rect 101426 426338 101662 426574
rect 101426 390658 101662 390894
rect 101426 390338 101662 390574
rect 101426 354658 101662 354894
rect 101426 354338 101662 354574
rect 101426 318658 101662 318894
rect 101426 318338 101662 318574
rect 101426 282658 101662 282894
rect 101426 282338 101662 282574
rect 101426 246658 101662 246894
rect 101426 246338 101662 246574
rect 101426 210658 101662 210894
rect 101426 210338 101662 210574
rect 101426 174658 101662 174894
rect 101426 174338 101662 174574
rect 101426 138658 101662 138894
rect 101426 138338 101662 138574
rect 101426 102658 101662 102894
rect 101426 102338 101662 102574
rect 101426 66658 101662 66894
rect 101426 66338 101662 66574
rect 101426 30658 101662 30894
rect 101426 30338 101662 30574
rect 83426 -6102 83662 -5866
rect 83426 -6422 83662 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112466 689698 112702 689934
rect 112466 689378 112702 689614
rect 112466 653698 112702 653934
rect 112466 653378 112702 653614
rect 112466 617698 112702 617934
rect 112466 617378 112702 617614
rect 112466 581698 112702 581934
rect 112466 581378 112702 581614
rect 112466 545698 112702 545934
rect 112466 545378 112702 545614
rect 112466 509698 112702 509934
rect 112466 509378 112702 509614
rect 112466 473698 112702 473934
rect 112466 473378 112702 473614
rect 112466 437698 112702 437934
rect 112466 437378 112702 437614
rect 112466 401698 112702 401934
rect 112466 401378 112702 401614
rect 112466 365698 112702 365934
rect 112466 365378 112702 365614
rect 112466 329698 112702 329934
rect 112466 329378 112702 329614
rect 112466 293698 112702 293934
rect 112466 293378 112702 293614
rect 112466 257698 112702 257934
rect 112466 257378 112702 257614
rect 112466 221698 112702 221934
rect 112466 221378 112702 221614
rect 112466 185698 112702 185934
rect 112466 185378 112702 185614
rect 112466 149698 112702 149934
rect 112466 149378 112702 149614
rect 112466 113698 112702 113934
rect 112466 113378 112702 113614
rect 112466 77698 112702 77934
rect 112466 77378 112702 77614
rect 112466 41698 112702 41934
rect 112466 41378 112702 41614
rect 112466 5698 112702 5934
rect 112466 5378 112702 5614
rect 112466 -2422 112702 -2186
rect 112466 -2742 112702 -2506
rect 115946 693178 116182 693414
rect 115946 692858 116182 693094
rect 115946 657178 116182 657414
rect 115946 656858 116182 657094
rect 115946 621178 116182 621414
rect 115946 620858 116182 621094
rect 115946 585178 116182 585414
rect 115946 584858 116182 585094
rect 115946 549178 116182 549414
rect 115946 548858 116182 549094
rect 115946 513178 116182 513414
rect 115946 512858 116182 513094
rect 115946 477178 116182 477414
rect 115946 476858 116182 477094
rect 115946 441178 116182 441414
rect 115946 440858 116182 441094
rect 115946 405178 116182 405414
rect 115946 404858 116182 405094
rect 115946 369178 116182 369414
rect 115946 368858 116182 369094
rect 115946 333178 116182 333414
rect 115946 332858 116182 333094
rect 115946 297178 116182 297414
rect 115946 296858 116182 297094
rect 115946 261178 116182 261414
rect 115946 260858 116182 261094
rect 115946 225178 116182 225414
rect 115946 224858 116182 225094
rect 115946 189178 116182 189414
rect 115946 188858 116182 189094
rect 115946 153178 116182 153414
rect 115946 152858 116182 153094
rect 115946 117178 116182 117414
rect 115946 116858 116182 117094
rect 115946 81178 116182 81414
rect 115946 80858 116182 81094
rect 115946 45178 116182 45414
rect 115946 44858 116182 45094
rect 115946 9178 116182 9414
rect 115946 8858 116182 9094
rect 115946 -4262 116182 -4026
rect 115946 -4582 116182 -4346
rect 137426 711042 137662 711278
rect 137426 710722 137662 710958
rect 133946 709202 134182 709438
rect 133946 708882 134182 709118
rect 130466 707362 130702 707598
rect 130466 707042 130702 707278
rect 119426 696658 119662 696894
rect 119426 696338 119662 696574
rect 119426 660658 119662 660894
rect 119426 660338 119662 660574
rect 119426 624658 119662 624894
rect 119426 624338 119662 624574
rect 119426 588658 119662 588894
rect 119426 588338 119662 588574
rect 119426 552658 119662 552894
rect 119426 552338 119662 552574
rect 119426 516658 119662 516894
rect 119426 516338 119662 516574
rect 119426 480658 119662 480894
rect 119426 480338 119662 480574
rect 119426 444658 119662 444894
rect 119426 444338 119662 444574
rect 119426 408658 119662 408894
rect 119426 408338 119662 408574
rect 119426 372658 119662 372894
rect 119426 372338 119662 372574
rect 119426 336658 119662 336894
rect 119426 336338 119662 336574
rect 119426 300658 119662 300894
rect 119426 300338 119662 300574
rect 119426 264658 119662 264894
rect 119426 264338 119662 264574
rect 119426 228658 119662 228894
rect 119426 228338 119662 228574
rect 119426 192658 119662 192894
rect 119426 192338 119662 192574
rect 119426 156658 119662 156894
rect 119426 156338 119662 156574
rect 119426 120658 119662 120894
rect 119426 120338 119662 120574
rect 119426 84658 119662 84894
rect 119426 84338 119662 84574
rect 119426 48658 119662 48894
rect 119426 48338 119662 48574
rect 119426 12658 119662 12894
rect 119426 12338 119662 12574
rect 101426 -7022 101662 -6786
rect 101426 -7342 101662 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130466 671698 130702 671934
rect 130466 671378 130702 671614
rect 130466 635698 130702 635934
rect 130466 635378 130702 635614
rect 130466 599698 130702 599934
rect 130466 599378 130702 599614
rect 130466 563698 130702 563934
rect 130466 563378 130702 563614
rect 130466 527698 130702 527934
rect 130466 527378 130702 527614
rect 130466 491698 130702 491934
rect 130466 491378 130702 491614
rect 130466 455698 130702 455934
rect 130466 455378 130702 455614
rect 130466 419698 130702 419934
rect 130466 419378 130702 419614
rect 130466 383698 130702 383934
rect 130466 383378 130702 383614
rect 130466 347698 130702 347934
rect 130466 347378 130702 347614
rect 130466 311698 130702 311934
rect 130466 311378 130702 311614
rect 130466 275698 130702 275934
rect 130466 275378 130702 275614
rect 130466 239698 130702 239934
rect 130466 239378 130702 239614
rect 130466 203698 130702 203934
rect 130466 203378 130702 203614
rect 130466 167698 130702 167934
rect 130466 167378 130702 167614
rect 130466 131698 130702 131934
rect 130466 131378 130702 131614
rect 130466 95698 130702 95934
rect 130466 95378 130702 95614
rect 130466 59698 130702 59934
rect 130466 59378 130702 59614
rect 130466 23698 130702 23934
rect 130466 23378 130702 23614
rect 130466 -3342 130702 -3106
rect 130466 -3662 130702 -3426
rect 133946 675178 134182 675414
rect 133946 674858 134182 675094
rect 133946 639178 134182 639414
rect 133946 638858 134182 639094
rect 133946 603178 134182 603414
rect 133946 602858 134182 603094
rect 133946 567178 134182 567414
rect 133946 566858 134182 567094
rect 133946 531178 134182 531414
rect 133946 530858 134182 531094
rect 133946 495178 134182 495414
rect 133946 494858 134182 495094
rect 133946 459178 134182 459414
rect 133946 458858 134182 459094
rect 133946 423178 134182 423414
rect 133946 422858 134182 423094
rect 133946 387178 134182 387414
rect 133946 386858 134182 387094
rect 133946 351178 134182 351414
rect 133946 350858 134182 351094
rect 133946 315178 134182 315414
rect 133946 314858 134182 315094
rect 133946 279178 134182 279414
rect 133946 278858 134182 279094
rect 133946 243178 134182 243414
rect 133946 242858 134182 243094
rect 133946 207178 134182 207414
rect 133946 206858 134182 207094
rect 133946 171178 134182 171414
rect 133946 170858 134182 171094
rect 133946 135178 134182 135414
rect 133946 134858 134182 135094
rect 133946 99178 134182 99414
rect 133946 98858 134182 99094
rect 133946 63178 134182 63414
rect 133946 62858 134182 63094
rect 133946 27178 134182 27414
rect 133946 26858 134182 27094
rect 133946 -5182 134182 -4946
rect 133946 -5502 134182 -5266
rect 155426 710122 155662 710358
rect 155426 709802 155662 710038
rect 151946 708282 152182 708518
rect 151946 707962 152182 708198
rect 148466 706442 148702 706678
rect 148466 706122 148702 706358
rect 137426 678658 137662 678894
rect 137426 678338 137662 678574
rect 137426 642658 137662 642894
rect 137426 642338 137662 642574
rect 137426 606658 137662 606894
rect 137426 606338 137662 606574
rect 137426 570658 137662 570894
rect 137426 570338 137662 570574
rect 137426 534658 137662 534894
rect 137426 534338 137662 534574
rect 137426 498658 137662 498894
rect 137426 498338 137662 498574
rect 137426 462658 137662 462894
rect 137426 462338 137662 462574
rect 137426 426658 137662 426894
rect 137426 426338 137662 426574
rect 137426 390658 137662 390894
rect 137426 390338 137662 390574
rect 137426 354658 137662 354894
rect 137426 354338 137662 354574
rect 137426 318658 137662 318894
rect 137426 318338 137662 318574
rect 137426 282658 137662 282894
rect 137426 282338 137662 282574
rect 137426 246658 137662 246894
rect 137426 246338 137662 246574
rect 137426 210658 137662 210894
rect 137426 210338 137662 210574
rect 137426 174658 137662 174894
rect 137426 174338 137662 174574
rect 137426 138658 137662 138894
rect 137426 138338 137662 138574
rect 137426 102658 137662 102894
rect 137426 102338 137662 102574
rect 137426 66658 137662 66894
rect 137426 66338 137662 66574
rect 137426 30658 137662 30894
rect 137426 30338 137662 30574
rect 119426 -6102 119662 -5866
rect 119426 -6422 119662 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148466 689698 148702 689934
rect 148466 689378 148702 689614
rect 148466 653698 148702 653934
rect 148466 653378 148702 653614
rect 148466 617698 148702 617934
rect 148466 617378 148702 617614
rect 148466 581698 148702 581934
rect 148466 581378 148702 581614
rect 148466 545698 148702 545934
rect 148466 545378 148702 545614
rect 148466 509698 148702 509934
rect 148466 509378 148702 509614
rect 148466 473698 148702 473934
rect 148466 473378 148702 473614
rect 148466 437698 148702 437934
rect 148466 437378 148702 437614
rect 148466 401698 148702 401934
rect 148466 401378 148702 401614
rect 148466 365698 148702 365934
rect 148466 365378 148702 365614
rect 148466 329698 148702 329934
rect 148466 329378 148702 329614
rect 148466 293698 148702 293934
rect 148466 293378 148702 293614
rect 148466 257698 148702 257934
rect 148466 257378 148702 257614
rect 148466 221698 148702 221934
rect 148466 221378 148702 221614
rect 148466 185698 148702 185934
rect 148466 185378 148702 185614
rect 148466 149698 148702 149934
rect 148466 149378 148702 149614
rect 148466 113698 148702 113934
rect 148466 113378 148702 113614
rect 148466 77698 148702 77934
rect 148466 77378 148702 77614
rect 148466 41698 148702 41934
rect 148466 41378 148702 41614
rect 148466 5698 148702 5934
rect 148466 5378 148702 5614
rect 148466 -2422 148702 -2186
rect 148466 -2742 148702 -2506
rect 151946 693178 152182 693414
rect 151946 692858 152182 693094
rect 151946 657178 152182 657414
rect 151946 656858 152182 657094
rect 151946 621178 152182 621414
rect 151946 620858 152182 621094
rect 151946 585178 152182 585414
rect 151946 584858 152182 585094
rect 151946 549178 152182 549414
rect 151946 548858 152182 549094
rect 151946 513178 152182 513414
rect 151946 512858 152182 513094
rect 151946 477178 152182 477414
rect 151946 476858 152182 477094
rect 151946 441178 152182 441414
rect 151946 440858 152182 441094
rect 151946 405178 152182 405414
rect 151946 404858 152182 405094
rect 151946 369178 152182 369414
rect 151946 368858 152182 369094
rect 151946 333178 152182 333414
rect 151946 332858 152182 333094
rect 151946 297178 152182 297414
rect 151946 296858 152182 297094
rect 151946 261178 152182 261414
rect 151946 260858 152182 261094
rect 151946 225178 152182 225414
rect 151946 224858 152182 225094
rect 151946 189178 152182 189414
rect 151946 188858 152182 189094
rect 151946 153178 152182 153414
rect 151946 152858 152182 153094
rect 151946 117178 152182 117414
rect 151946 116858 152182 117094
rect 151946 81178 152182 81414
rect 151946 80858 152182 81094
rect 151946 45178 152182 45414
rect 151946 44858 152182 45094
rect 151946 9178 152182 9414
rect 151946 8858 152182 9094
rect 151946 -4262 152182 -4026
rect 151946 -4582 152182 -4346
rect 173426 711042 173662 711278
rect 173426 710722 173662 710958
rect 169946 709202 170182 709438
rect 169946 708882 170182 709118
rect 166466 707362 166702 707598
rect 166466 707042 166702 707278
rect 155426 696658 155662 696894
rect 155426 696338 155662 696574
rect 155426 660658 155662 660894
rect 155426 660338 155662 660574
rect 155426 624658 155662 624894
rect 155426 624338 155662 624574
rect 155426 588658 155662 588894
rect 155426 588338 155662 588574
rect 155426 552658 155662 552894
rect 155426 552338 155662 552574
rect 155426 516658 155662 516894
rect 155426 516338 155662 516574
rect 155426 480658 155662 480894
rect 155426 480338 155662 480574
rect 155426 444658 155662 444894
rect 155426 444338 155662 444574
rect 155426 408658 155662 408894
rect 155426 408338 155662 408574
rect 155426 372658 155662 372894
rect 155426 372338 155662 372574
rect 155426 336658 155662 336894
rect 155426 336338 155662 336574
rect 155426 300658 155662 300894
rect 155426 300338 155662 300574
rect 155426 264658 155662 264894
rect 155426 264338 155662 264574
rect 155426 228658 155662 228894
rect 155426 228338 155662 228574
rect 155426 192658 155662 192894
rect 155426 192338 155662 192574
rect 155426 156658 155662 156894
rect 155426 156338 155662 156574
rect 155426 120658 155662 120894
rect 155426 120338 155662 120574
rect 155426 84658 155662 84894
rect 155426 84338 155662 84574
rect 155426 48658 155662 48894
rect 155426 48338 155662 48574
rect 155426 12658 155662 12894
rect 155426 12338 155662 12574
rect 137426 -7022 137662 -6786
rect 137426 -7342 137662 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166466 671698 166702 671934
rect 166466 671378 166702 671614
rect 166466 635698 166702 635934
rect 166466 635378 166702 635614
rect 166466 599698 166702 599934
rect 166466 599378 166702 599614
rect 166466 563698 166702 563934
rect 166466 563378 166702 563614
rect 166466 527698 166702 527934
rect 166466 527378 166702 527614
rect 166466 491698 166702 491934
rect 166466 491378 166702 491614
rect 166466 455698 166702 455934
rect 166466 455378 166702 455614
rect 166466 419698 166702 419934
rect 166466 419378 166702 419614
rect 166466 383698 166702 383934
rect 166466 383378 166702 383614
rect 166466 347698 166702 347934
rect 166466 347378 166702 347614
rect 166466 311698 166702 311934
rect 166466 311378 166702 311614
rect 166466 275698 166702 275934
rect 166466 275378 166702 275614
rect 166466 239698 166702 239934
rect 166466 239378 166702 239614
rect 166466 203698 166702 203934
rect 166466 203378 166702 203614
rect 166466 167698 166702 167934
rect 166466 167378 166702 167614
rect 166466 131698 166702 131934
rect 166466 131378 166702 131614
rect 166466 95698 166702 95934
rect 166466 95378 166702 95614
rect 166466 59698 166702 59934
rect 166466 59378 166702 59614
rect 166466 23698 166702 23934
rect 166466 23378 166702 23614
rect 166466 -3342 166702 -3106
rect 166466 -3662 166702 -3426
rect 169946 675178 170182 675414
rect 169946 674858 170182 675094
rect 169946 639178 170182 639414
rect 169946 638858 170182 639094
rect 169946 603178 170182 603414
rect 169946 602858 170182 603094
rect 169946 567178 170182 567414
rect 169946 566858 170182 567094
rect 169946 531178 170182 531414
rect 169946 530858 170182 531094
rect 169946 495178 170182 495414
rect 169946 494858 170182 495094
rect 169946 459178 170182 459414
rect 169946 458858 170182 459094
rect 169946 423178 170182 423414
rect 169946 422858 170182 423094
rect 169946 387178 170182 387414
rect 169946 386858 170182 387094
rect 169946 351178 170182 351414
rect 169946 350858 170182 351094
rect 169946 315178 170182 315414
rect 169946 314858 170182 315094
rect 169946 279178 170182 279414
rect 169946 278858 170182 279094
rect 169946 243178 170182 243414
rect 169946 242858 170182 243094
rect 169946 207178 170182 207414
rect 169946 206858 170182 207094
rect 169946 171178 170182 171414
rect 169946 170858 170182 171094
rect 169946 135178 170182 135414
rect 169946 134858 170182 135094
rect 169946 99178 170182 99414
rect 169946 98858 170182 99094
rect 169946 63178 170182 63414
rect 169946 62858 170182 63094
rect 169946 27178 170182 27414
rect 169946 26858 170182 27094
rect 169946 -5182 170182 -4946
rect 169946 -5502 170182 -5266
rect 191426 710122 191662 710358
rect 191426 709802 191662 710038
rect 187946 708282 188182 708518
rect 187946 707962 188182 708198
rect 184466 706442 184702 706678
rect 184466 706122 184702 706358
rect 173426 678658 173662 678894
rect 173426 678338 173662 678574
rect 173426 642658 173662 642894
rect 173426 642338 173662 642574
rect 173426 606658 173662 606894
rect 173426 606338 173662 606574
rect 173426 570658 173662 570894
rect 173426 570338 173662 570574
rect 173426 534658 173662 534894
rect 173426 534338 173662 534574
rect 173426 498658 173662 498894
rect 173426 498338 173662 498574
rect 173426 462658 173662 462894
rect 173426 462338 173662 462574
rect 173426 426658 173662 426894
rect 173426 426338 173662 426574
rect 173426 390658 173662 390894
rect 173426 390338 173662 390574
rect 173426 354658 173662 354894
rect 173426 354338 173662 354574
rect 173426 318658 173662 318894
rect 173426 318338 173662 318574
rect 173426 282658 173662 282894
rect 173426 282338 173662 282574
rect 173426 246658 173662 246894
rect 173426 246338 173662 246574
rect 173426 210658 173662 210894
rect 173426 210338 173662 210574
rect 173426 174658 173662 174894
rect 173426 174338 173662 174574
rect 173426 138658 173662 138894
rect 173426 138338 173662 138574
rect 173426 102658 173662 102894
rect 173426 102338 173662 102574
rect 173426 66658 173662 66894
rect 173426 66338 173662 66574
rect 173426 30658 173662 30894
rect 173426 30338 173662 30574
rect 155426 -6102 155662 -5866
rect 155426 -6422 155662 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184466 689698 184702 689934
rect 184466 689378 184702 689614
rect 184466 653698 184702 653934
rect 184466 653378 184702 653614
rect 184466 617698 184702 617934
rect 184466 617378 184702 617614
rect 184466 581698 184702 581934
rect 184466 581378 184702 581614
rect 184466 545698 184702 545934
rect 184466 545378 184702 545614
rect 184466 509698 184702 509934
rect 184466 509378 184702 509614
rect 184466 473698 184702 473934
rect 184466 473378 184702 473614
rect 184466 437698 184702 437934
rect 184466 437378 184702 437614
rect 184466 401698 184702 401934
rect 184466 401378 184702 401614
rect 184466 365698 184702 365934
rect 184466 365378 184702 365614
rect 184466 329698 184702 329934
rect 184466 329378 184702 329614
rect 184466 293698 184702 293934
rect 184466 293378 184702 293614
rect 184466 257698 184702 257934
rect 184466 257378 184702 257614
rect 184466 221698 184702 221934
rect 184466 221378 184702 221614
rect 184466 185698 184702 185934
rect 184466 185378 184702 185614
rect 184466 149698 184702 149934
rect 184466 149378 184702 149614
rect 184466 113698 184702 113934
rect 184466 113378 184702 113614
rect 184466 77698 184702 77934
rect 184466 77378 184702 77614
rect 184466 41698 184702 41934
rect 184466 41378 184702 41614
rect 184466 5698 184702 5934
rect 184466 5378 184702 5614
rect 184466 -2422 184702 -2186
rect 184466 -2742 184702 -2506
rect 187946 693178 188182 693414
rect 187946 692858 188182 693094
rect 187946 657178 188182 657414
rect 187946 656858 188182 657094
rect 187946 621178 188182 621414
rect 187946 620858 188182 621094
rect 187946 585178 188182 585414
rect 187946 584858 188182 585094
rect 187946 549178 188182 549414
rect 187946 548858 188182 549094
rect 187946 513178 188182 513414
rect 187946 512858 188182 513094
rect 187946 477178 188182 477414
rect 187946 476858 188182 477094
rect 187946 441178 188182 441414
rect 187946 440858 188182 441094
rect 187946 405178 188182 405414
rect 187946 404858 188182 405094
rect 187946 369178 188182 369414
rect 187946 368858 188182 369094
rect 187946 333178 188182 333414
rect 187946 332858 188182 333094
rect 187946 297178 188182 297414
rect 187946 296858 188182 297094
rect 187946 261178 188182 261414
rect 187946 260858 188182 261094
rect 187946 225178 188182 225414
rect 187946 224858 188182 225094
rect 187946 189178 188182 189414
rect 187946 188858 188182 189094
rect 187946 153178 188182 153414
rect 187946 152858 188182 153094
rect 187946 117178 188182 117414
rect 187946 116858 188182 117094
rect 187946 81178 188182 81414
rect 187946 80858 188182 81094
rect 187946 45178 188182 45414
rect 187946 44858 188182 45094
rect 187946 9178 188182 9414
rect 187946 8858 188182 9094
rect 187946 -4262 188182 -4026
rect 187946 -4582 188182 -4346
rect 209426 711042 209662 711278
rect 209426 710722 209662 710958
rect 205946 709202 206182 709438
rect 205946 708882 206182 709118
rect 202466 707362 202702 707598
rect 202466 707042 202702 707278
rect 191426 696658 191662 696894
rect 191426 696338 191662 696574
rect 191426 660658 191662 660894
rect 191426 660338 191662 660574
rect 191426 624658 191662 624894
rect 191426 624338 191662 624574
rect 191426 588658 191662 588894
rect 191426 588338 191662 588574
rect 191426 552658 191662 552894
rect 191426 552338 191662 552574
rect 191426 516658 191662 516894
rect 191426 516338 191662 516574
rect 191426 480658 191662 480894
rect 191426 480338 191662 480574
rect 191426 444658 191662 444894
rect 191426 444338 191662 444574
rect 191426 408658 191662 408894
rect 191426 408338 191662 408574
rect 191426 372658 191662 372894
rect 191426 372338 191662 372574
rect 191426 336658 191662 336894
rect 191426 336338 191662 336574
rect 191426 300658 191662 300894
rect 191426 300338 191662 300574
rect 191426 264658 191662 264894
rect 191426 264338 191662 264574
rect 191426 228658 191662 228894
rect 191426 228338 191662 228574
rect 191426 192658 191662 192894
rect 191426 192338 191662 192574
rect 191426 156658 191662 156894
rect 191426 156338 191662 156574
rect 191426 120658 191662 120894
rect 191426 120338 191662 120574
rect 191426 84658 191662 84894
rect 191426 84338 191662 84574
rect 191426 48658 191662 48894
rect 191426 48338 191662 48574
rect 191426 12658 191662 12894
rect 191426 12338 191662 12574
rect 173426 -7022 173662 -6786
rect 173426 -7342 173662 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202466 671698 202702 671934
rect 202466 671378 202702 671614
rect 202466 635698 202702 635934
rect 202466 635378 202702 635614
rect 202466 599698 202702 599934
rect 202466 599378 202702 599614
rect 202466 563698 202702 563934
rect 202466 563378 202702 563614
rect 202466 527698 202702 527934
rect 202466 527378 202702 527614
rect 202466 491698 202702 491934
rect 202466 491378 202702 491614
rect 202466 455698 202702 455934
rect 202466 455378 202702 455614
rect 202466 419698 202702 419934
rect 202466 419378 202702 419614
rect 202466 383698 202702 383934
rect 202466 383378 202702 383614
rect 202466 347698 202702 347934
rect 202466 347378 202702 347614
rect 202466 311698 202702 311934
rect 202466 311378 202702 311614
rect 202466 275698 202702 275934
rect 202466 275378 202702 275614
rect 202466 239698 202702 239934
rect 202466 239378 202702 239614
rect 202466 203698 202702 203934
rect 202466 203378 202702 203614
rect 202466 167698 202702 167934
rect 202466 167378 202702 167614
rect 202466 131698 202702 131934
rect 202466 131378 202702 131614
rect 202466 95698 202702 95934
rect 202466 95378 202702 95614
rect 202466 59698 202702 59934
rect 202466 59378 202702 59614
rect 202466 23698 202702 23934
rect 202466 23378 202702 23614
rect 202466 -3342 202702 -3106
rect 202466 -3662 202702 -3426
rect 205946 675178 206182 675414
rect 205946 674858 206182 675094
rect 205946 639178 206182 639414
rect 205946 638858 206182 639094
rect 205946 603178 206182 603414
rect 205946 602858 206182 603094
rect 205946 567178 206182 567414
rect 205946 566858 206182 567094
rect 205946 531178 206182 531414
rect 205946 530858 206182 531094
rect 205946 495178 206182 495414
rect 205946 494858 206182 495094
rect 205946 459178 206182 459414
rect 205946 458858 206182 459094
rect 205946 423178 206182 423414
rect 205946 422858 206182 423094
rect 205946 387178 206182 387414
rect 205946 386858 206182 387094
rect 205946 351178 206182 351414
rect 205946 350858 206182 351094
rect 205946 315178 206182 315414
rect 205946 314858 206182 315094
rect 205946 279178 206182 279414
rect 205946 278858 206182 279094
rect 205946 243178 206182 243414
rect 205946 242858 206182 243094
rect 205946 207178 206182 207414
rect 205946 206858 206182 207094
rect 205946 171178 206182 171414
rect 205946 170858 206182 171094
rect 205946 135178 206182 135414
rect 205946 134858 206182 135094
rect 205946 99178 206182 99414
rect 205946 98858 206182 99094
rect 205946 63178 206182 63414
rect 205946 62858 206182 63094
rect 205946 27178 206182 27414
rect 205946 26858 206182 27094
rect 205946 -5182 206182 -4946
rect 205946 -5502 206182 -5266
rect 227426 710122 227662 710358
rect 227426 709802 227662 710038
rect 223946 708282 224182 708518
rect 223946 707962 224182 708198
rect 220466 706442 220702 706678
rect 220466 706122 220702 706358
rect 209426 678658 209662 678894
rect 209426 678338 209662 678574
rect 209426 642658 209662 642894
rect 209426 642338 209662 642574
rect 209426 606658 209662 606894
rect 209426 606338 209662 606574
rect 209426 570658 209662 570894
rect 209426 570338 209662 570574
rect 209426 534658 209662 534894
rect 209426 534338 209662 534574
rect 209426 498658 209662 498894
rect 209426 498338 209662 498574
rect 209426 462658 209662 462894
rect 209426 462338 209662 462574
rect 209426 426658 209662 426894
rect 209426 426338 209662 426574
rect 209426 390658 209662 390894
rect 209426 390338 209662 390574
rect 209426 354658 209662 354894
rect 209426 354338 209662 354574
rect 209426 318658 209662 318894
rect 209426 318338 209662 318574
rect 209426 282658 209662 282894
rect 209426 282338 209662 282574
rect 209426 246658 209662 246894
rect 209426 246338 209662 246574
rect 209426 210658 209662 210894
rect 209426 210338 209662 210574
rect 209426 174658 209662 174894
rect 209426 174338 209662 174574
rect 209426 138658 209662 138894
rect 209426 138338 209662 138574
rect 209426 102658 209662 102894
rect 209426 102338 209662 102574
rect 209426 66658 209662 66894
rect 209426 66338 209662 66574
rect 209426 30658 209662 30894
rect 209426 30338 209662 30574
rect 191426 -6102 191662 -5866
rect 191426 -6422 191662 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220466 689698 220702 689934
rect 220466 689378 220702 689614
rect 220466 653698 220702 653934
rect 220466 653378 220702 653614
rect 220466 617698 220702 617934
rect 220466 617378 220702 617614
rect 220466 581698 220702 581934
rect 220466 581378 220702 581614
rect 220466 545698 220702 545934
rect 220466 545378 220702 545614
rect 220466 509698 220702 509934
rect 220466 509378 220702 509614
rect 220466 473698 220702 473934
rect 220466 473378 220702 473614
rect 220466 437698 220702 437934
rect 220466 437378 220702 437614
rect 220466 401698 220702 401934
rect 220466 401378 220702 401614
rect 220466 365698 220702 365934
rect 220466 365378 220702 365614
rect 220466 329698 220702 329934
rect 220466 329378 220702 329614
rect 220466 293698 220702 293934
rect 220466 293378 220702 293614
rect 220466 257698 220702 257934
rect 220466 257378 220702 257614
rect 220466 221698 220702 221934
rect 220466 221378 220702 221614
rect 220466 185698 220702 185934
rect 220466 185378 220702 185614
rect 220466 149698 220702 149934
rect 220466 149378 220702 149614
rect 220466 113698 220702 113934
rect 220466 113378 220702 113614
rect 220466 77698 220702 77934
rect 220466 77378 220702 77614
rect 220466 41698 220702 41934
rect 220466 41378 220702 41614
rect 220466 5698 220702 5934
rect 220466 5378 220702 5614
rect 220466 -2422 220702 -2186
rect 220466 -2742 220702 -2506
rect 223946 693178 224182 693414
rect 223946 692858 224182 693094
rect 223946 657178 224182 657414
rect 223946 656858 224182 657094
rect 223946 621178 224182 621414
rect 223946 620858 224182 621094
rect 223946 585178 224182 585414
rect 223946 584858 224182 585094
rect 223946 549178 224182 549414
rect 223946 548858 224182 549094
rect 223946 513178 224182 513414
rect 223946 512858 224182 513094
rect 223946 477178 224182 477414
rect 223946 476858 224182 477094
rect 223946 441178 224182 441414
rect 223946 440858 224182 441094
rect 223946 405178 224182 405414
rect 223946 404858 224182 405094
rect 223946 369178 224182 369414
rect 223946 368858 224182 369094
rect 223946 333178 224182 333414
rect 223946 332858 224182 333094
rect 223946 297178 224182 297414
rect 223946 296858 224182 297094
rect 223946 261178 224182 261414
rect 223946 260858 224182 261094
rect 223946 225178 224182 225414
rect 223946 224858 224182 225094
rect 223946 189178 224182 189414
rect 223946 188858 224182 189094
rect 223946 153178 224182 153414
rect 223946 152858 224182 153094
rect 223946 117178 224182 117414
rect 223946 116858 224182 117094
rect 223946 81178 224182 81414
rect 223946 80858 224182 81094
rect 223946 45178 224182 45414
rect 223946 44858 224182 45094
rect 223946 9178 224182 9414
rect 223946 8858 224182 9094
rect 223946 -4262 224182 -4026
rect 223946 -4582 224182 -4346
rect 245426 711042 245662 711278
rect 245426 710722 245662 710958
rect 241946 709202 242182 709438
rect 241946 708882 242182 709118
rect 238466 707362 238702 707598
rect 238466 707042 238702 707278
rect 227426 696658 227662 696894
rect 227426 696338 227662 696574
rect 227426 660658 227662 660894
rect 227426 660338 227662 660574
rect 227426 624658 227662 624894
rect 227426 624338 227662 624574
rect 227426 588658 227662 588894
rect 227426 588338 227662 588574
rect 227426 552658 227662 552894
rect 227426 552338 227662 552574
rect 227426 516658 227662 516894
rect 227426 516338 227662 516574
rect 227426 480658 227662 480894
rect 227426 480338 227662 480574
rect 227426 444658 227662 444894
rect 227426 444338 227662 444574
rect 227426 408658 227662 408894
rect 227426 408338 227662 408574
rect 227426 372658 227662 372894
rect 227426 372338 227662 372574
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 230710 360622 230946 360858
rect 227426 336658 227662 336894
rect 227426 336338 227662 336574
rect 227426 300658 227662 300894
rect 227426 300338 227662 300574
rect 227426 264658 227662 264894
rect 227426 264338 227662 264574
rect 227426 228658 227662 228894
rect 227426 228338 227662 228574
rect 227426 192658 227662 192894
rect 227426 192338 227662 192574
rect 227426 156658 227662 156894
rect 227426 156338 227662 156574
rect 227426 120658 227662 120894
rect 227426 120338 227662 120574
rect 227426 84658 227662 84894
rect 227426 84338 227662 84574
rect 227426 48658 227662 48894
rect 227426 48338 227662 48574
rect 227426 12658 227662 12894
rect 227426 12338 227662 12574
rect 209426 -7022 209662 -6786
rect 209426 -7342 209662 -7106
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238466 671698 238702 671934
rect 238466 671378 238702 671614
rect 238466 635698 238702 635934
rect 238466 635378 238702 635614
rect 238466 599698 238702 599934
rect 238466 599378 238702 599614
rect 238466 563698 238702 563934
rect 238466 563378 238702 563614
rect 238466 527698 238702 527934
rect 238466 527378 238702 527614
rect 238466 491698 238702 491934
rect 238466 491378 238702 491614
rect 238466 455698 238702 455934
rect 238466 455378 238702 455614
rect 238466 419698 238702 419934
rect 238466 419378 238702 419614
rect 238466 383698 238702 383934
rect 238466 383378 238702 383614
rect 241946 675178 242182 675414
rect 241946 674858 242182 675094
rect 241946 639178 242182 639414
rect 241946 638858 242182 639094
rect 241946 603178 242182 603414
rect 241946 602858 242182 603094
rect 241946 567178 242182 567414
rect 241946 566858 242182 567094
rect 241946 531178 242182 531414
rect 241946 530858 242182 531094
rect 241946 495178 242182 495414
rect 241946 494858 242182 495094
rect 241946 459178 242182 459414
rect 241946 458858 242182 459094
rect 241946 423178 242182 423414
rect 241946 422858 242182 423094
rect 241946 387178 242182 387414
rect 241946 386858 242182 387094
rect 238990 363342 239226 363578
rect 238990 360622 239226 360858
rect 238466 347698 238702 347934
rect 238466 347378 238702 347614
rect 238466 311698 238702 311934
rect 238466 311378 238702 311614
rect 238466 275698 238702 275934
rect 238466 275378 238702 275614
rect 238466 239698 238702 239934
rect 238466 239378 238702 239614
rect 238466 203698 238702 203934
rect 238466 203378 238702 203614
rect 238466 167698 238702 167934
rect 238466 167378 238702 167614
rect 238466 131698 238702 131934
rect 238466 131378 238702 131614
rect 238466 95698 238702 95934
rect 238466 95378 238702 95614
rect 238466 59698 238702 59934
rect 238466 59378 238702 59614
rect 238466 23698 238702 23934
rect 238466 23378 238702 23614
rect 238466 -3342 238702 -3106
rect 238466 -3662 238702 -3426
rect 241946 351178 242182 351414
rect 241946 350858 242182 351094
rect 241946 315178 242182 315414
rect 241946 314858 242182 315094
rect 241946 279178 242182 279414
rect 241946 278858 242182 279094
rect 241946 243178 242182 243414
rect 241946 242858 242182 243094
rect 241946 207178 242182 207414
rect 241946 206858 242182 207094
rect 241946 171178 242182 171414
rect 241946 170858 242182 171094
rect 241946 135178 242182 135414
rect 241946 134858 242182 135094
rect 241946 99178 242182 99414
rect 241946 98858 242182 99094
rect 241946 63178 242182 63414
rect 241946 62858 242182 63094
rect 241946 27178 242182 27414
rect 241946 26858 242182 27094
rect 241946 -5182 242182 -4946
rect 241946 -5502 242182 -5266
rect 263426 710122 263662 710358
rect 263426 709802 263662 710038
rect 259946 708282 260182 708518
rect 259946 707962 260182 708198
rect 256466 706442 256702 706678
rect 256466 706122 256702 706358
rect 245426 678658 245662 678894
rect 245426 678338 245662 678574
rect 245426 642658 245662 642894
rect 245426 642338 245662 642574
rect 245426 606658 245662 606894
rect 245426 606338 245662 606574
rect 245426 570658 245662 570894
rect 245426 570338 245662 570574
rect 245426 534658 245662 534894
rect 245426 534338 245662 534574
rect 245426 498658 245662 498894
rect 245426 498338 245662 498574
rect 245426 462658 245662 462894
rect 245426 462338 245662 462574
rect 245426 426658 245662 426894
rect 245426 426338 245662 426574
rect 245426 390658 245662 390894
rect 245426 390338 245662 390574
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 248558 363342 248794 363578
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 248558 360622 248794 360858
rect 245426 354658 245662 354894
rect 245426 354338 245662 354574
rect 245426 318658 245662 318894
rect 245426 318338 245662 318574
rect 245426 282658 245662 282894
rect 245426 282338 245662 282574
rect 245426 246658 245662 246894
rect 245426 246338 245662 246574
rect 245426 210658 245662 210894
rect 245426 210338 245662 210574
rect 245426 174658 245662 174894
rect 245426 174338 245662 174574
rect 245426 138658 245662 138894
rect 245426 138338 245662 138574
rect 245426 102658 245662 102894
rect 245426 102338 245662 102574
rect 245426 66658 245662 66894
rect 245426 66338 245662 66574
rect 245426 30658 245662 30894
rect 245426 30338 245662 30574
rect 227426 -6102 227662 -5866
rect 227426 -6422 227662 -6186
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256466 689698 256702 689934
rect 256466 689378 256702 689614
rect 256466 653698 256702 653934
rect 256466 653378 256702 653614
rect 256466 617698 256702 617934
rect 256466 617378 256702 617614
rect 256466 581698 256702 581934
rect 256466 581378 256702 581614
rect 256466 545698 256702 545934
rect 256466 545378 256702 545614
rect 256466 509698 256702 509934
rect 256466 509378 256702 509614
rect 256466 473698 256702 473934
rect 256466 473378 256702 473614
rect 256466 437698 256702 437934
rect 256466 437378 256702 437614
rect 256466 401698 256702 401934
rect 256466 401378 256702 401614
rect 256466 365698 256702 365934
rect 256466 365378 256702 365614
rect 256466 329698 256702 329934
rect 256466 329378 256702 329614
rect 256466 293698 256702 293934
rect 256466 293378 256702 293614
rect 256466 257698 256702 257934
rect 256466 257378 256702 257614
rect 256466 221698 256702 221934
rect 256466 221378 256702 221614
rect 256466 185698 256702 185934
rect 256466 185378 256702 185614
rect 256466 149698 256702 149934
rect 256466 149378 256702 149614
rect 256466 113698 256702 113934
rect 256466 113378 256702 113614
rect 256466 77698 256702 77934
rect 256466 77378 256702 77614
rect 256466 41698 256702 41934
rect 256466 41378 256702 41614
rect 256466 5698 256702 5934
rect 256466 5378 256702 5614
rect 256466 -2422 256702 -2186
rect 256466 -2742 256702 -2506
rect 259946 693178 260182 693414
rect 259946 692858 260182 693094
rect 259946 657178 260182 657414
rect 259946 656858 260182 657094
rect 259946 621178 260182 621414
rect 259946 620858 260182 621094
rect 259946 585178 260182 585414
rect 259946 584858 260182 585094
rect 259946 549178 260182 549414
rect 259946 548858 260182 549094
rect 259946 513178 260182 513414
rect 259946 512858 260182 513094
rect 259946 477178 260182 477414
rect 259946 476858 260182 477094
rect 259946 441178 260182 441414
rect 259946 440858 260182 441094
rect 259946 405178 260182 405414
rect 259946 404858 260182 405094
rect 259946 369178 260182 369414
rect 259946 368858 260182 369094
rect 259946 333178 260182 333414
rect 259946 332858 260182 333094
rect 259946 297178 260182 297414
rect 259946 296858 260182 297094
rect 259946 261178 260182 261414
rect 259946 260858 260182 261094
rect 259946 225178 260182 225414
rect 259946 224858 260182 225094
rect 259946 189178 260182 189414
rect 259946 188858 260182 189094
rect 259946 153178 260182 153414
rect 259946 152858 260182 153094
rect 259946 117178 260182 117414
rect 259946 116858 260182 117094
rect 259946 81178 260182 81414
rect 259946 80858 260182 81094
rect 259946 45178 260182 45414
rect 259946 44858 260182 45094
rect 259946 9178 260182 9414
rect 259946 8858 260182 9094
rect 259946 -4262 260182 -4026
rect 259946 -4582 260182 -4346
rect 281426 711042 281662 711278
rect 281426 710722 281662 710958
rect 277946 709202 278182 709438
rect 277946 708882 278182 709118
rect 274466 707362 274702 707598
rect 274466 707042 274702 707278
rect 263426 696658 263662 696894
rect 263426 696338 263662 696574
rect 263426 660658 263662 660894
rect 263426 660338 263662 660574
rect 263426 624658 263662 624894
rect 263426 624338 263662 624574
rect 263426 588658 263662 588894
rect 263426 588338 263662 588574
rect 263426 552658 263662 552894
rect 263426 552338 263662 552574
rect 263426 516658 263662 516894
rect 263426 516338 263662 516574
rect 263426 480658 263662 480894
rect 263426 480338 263662 480574
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 263426 444658 263662 444894
rect 263426 444338 263662 444574
rect 263426 408658 263662 408894
rect 263426 408338 263662 408574
rect 263426 372658 263662 372894
rect 263426 372338 263662 372574
rect 263426 336658 263662 336894
rect 263426 336338 263662 336574
rect 263426 300658 263662 300894
rect 263426 300338 263662 300574
rect 263426 264658 263662 264894
rect 263426 264338 263662 264574
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 268798 363342 269034 363578
rect 268798 360622 269034 360858
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 263426 228658 263662 228894
rect 263426 228338 263662 228574
rect 263426 192658 263662 192894
rect 263426 192338 263662 192574
rect 263426 156658 263662 156894
rect 263426 156338 263662 156574
rect 263426 120658 263662 120894
rect 263426 120338 263662 120574
rect 263426 84658 263662 84894
rect 263426 84338 263662 84574
rect 263426 48658 263662 48894
rect 263426 48338 263662 48574
rect 263426 12658 263662 12894
rect 263426 12338 263662 12574
rect 245426 -7022 245662 -6786
rect 245426 -7342 245662 -7106
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274466 671698 274702 671934
rect 274466 671378 274702 671614
rect 274466 635698 274702 635934
rect 274466 635378 274702 635614
rect 274466 599698 274702 599934
rect 274466 599378 274702 599614
rect 274466 563698 274702 563934
rect 274466 563378 274702 563614
rect 274466 527698 274702 527934
rect 274466 527378 274702 527614
rect 274466 491698 274702 491934
rect 274466 491378 274702 491614
rect 274466 455698 274702 455934
rect 274466 455378 274702 455614
rect 274466 419698 274702 419934
rect 274466 419378 274702 419614
rect 274466 383698 274702 383934
rect 274466 383378 274702 383614
rect 274466 347698 274702 347934
rect 274466 347378 274702 347614
rect 274466 311698 274702 311934
rect 274466 311378 274702 311614
rect 274466 275698 274702 275934
rect 274466 275378 274702 275614
rect 274466 239698 274702 239934
rect 274466 239378 274702 239614
rect 274466 203698 274702 203934
rect 274466 203378 274702 203614
rect 274466 167698 274702 167934
rect 274466 167378 274702 167614
rect 274466 131698 274702 131934
rect 274466 131378 274702 131614
rect 274466 95698 274702 95934
rect 274466 95378 274702 95614
rect 274466 59698 274702 59934
rect 274466 59378 274702 59614
rect 274466 23698 274702 23934
rect 274466 23378 274702 23614
rect 274466 -3342 274702 -3106
rect 274466 -3662 274702 -3426
rect 277946 675178 278182 675414
rect 277946 674858 278182 675094
rect 277946 639178 278182 639414
rect 277946 638858 278182 639094
rect 277946 603178 278182 603414
rect 277946 602858 278182 603094
rect 277946 567178 278182 567414
rect 277946 566858 278182 567094
rect 277946 531178 278182 531414
rect 277946 530858 278182 531094
rect 277946 495178 278182 495414
rect 277946 494858 278182 495094
rect 277946 459178 278182 459414
rect 277946 458858 278182 459094
rect 277946 423178 278182 423414
rect 277946 422858 278182 423094
rect 277946 387178 278182 387414
rect 277946 386858 278182 387094
rect 277946 351178 278182 351414
rect 277946 350858 278182 351094
rect 277946 315178 278182 315414
rect 277946 314858 278182 315094
rect 277946 279178 278182 279414
rect 277946 278858 278182 279094
rect 277946 243178 278182 243414
rect 277946 242858 278182 243094
rect 277946 207178 278182 207414
rect 277946 206858 278182 207094
rect 277946 171178 278182 171414
rect 277946 170858 278182 171094
rect 277946 135178 278182 135414
rect 277946 134858 278182 135094
rect 277946 99178 278182 99414
rect 277946 98858 278182 99094
rect 277946 63178 278182 63414
rect 277946 62858 278182 63094
rect 277946 27178 278182 27414
rect 277946 26858 278182 27094
rect 277946 -5182 278182 -4946
rect 277946 -5502 278182 -5266
rect 299426 710122 299662 710358
rect 299426 709802 299662 710038
rect 295946 708282 296182 708518
rect 295946 707962 296182 708198
rect 292466 706442 292702 706678
rect 292466 706122 292702 706358
rect 281426 678658 281662 678894
rect 281426 678338 281662 678574
rect 281426 642658 281662 642894
rect 281426 642338 281662 642574
rect 281426 606658 281662 606894
rect 281426 606338 281662 606574
rect 281426 570658 281662 570894
rect 281426 570338 281662 570574
rect 281426 534658 281662 534894
rect 281426 534338 281662 534574
rect 281426 498658 281662 498894
rect 281426 498338 281662 498574
rect 281426 462658 281662 462894
rect 281426 462338 281662 462574
rect 281426 426658 281662 426894
rect 281426 426338 281662 426574
rect 281426 390658 281662 390894
rect 281426 390338 281662 390574
rect 281426 354658 281662 354894
rect 281426 354338 281662 354574
rect 281426 318658 281662 318894
rect 281426 318338 281662 318574
rect 281426 282658 281662 282894
rect 281426 282338 281662 282574
rect 281426 246658 281662 246894
rect 281426 246338 281662 246574
rect 281426 210658 281662 210894
rect 281426 210338 281662 210574
rect 281426 174658 281662 174894
rect 281426 174338 281662 174574
rect 281426 138658 281662 138894
rect 281426 138338 281662 138574
rect 281426 102658 281662 102894
rect 281426 102338 281662 102574
rect 281426 66658 281662 66894
rect 281426 66338 281662 66574
rect 281426 30658 281662 30894
rect 281426 30338 281662 30574
rect 263426 -6102 263662 -5866
rect 263426 -6422 263662 -6186
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292466 689698 292702 689934
rect 292466 689378 292702 689614
rect 292466 653698 292702 653934
rect 292466 653378 292702 653614
rect 292466 617698 292702 617934
rect 292466 617378 292702 617614
rect 292466 581698 292702 581934
rect 292466 581378 292702 581614
rect 292466 545698 292702 545934
rect 292466 545378 292702 545614
rect 292466 509698 292702 509934
rect 292466 509378 292702 509614
rect 292466 473698 292702 473934
rect 292466 473378 292702 473614
rect 292466 437698 292702 437934
rect 292466 437378 292702 437614
rect 292466 401698 292702 401934
rect 292466 401378 292702 401614
rect 292466 365698 292702 365934
rect 292466 365378 292702 365614
rect 292466 329698 292702 329934
rect 292466 329378 292702 329614
rect 292466 293698 292702 293934
rect 292466 293378 292702 293614
rect 292466 257698 292702 257934
rect 292466 257378 292702 257614
rect 292466 221698 292702 221934
rect 292466 221378 292702 221614
rect 292466 185698 292702 185934
rect 292466 185378 292702 185614
rect 292466 149698 292702 149934
rect 292466 149378 292702 149614
rect 292466 113698 292702 113934
rect 292466 113378 292702 113614
rect 292466 77698 292702 77934
rect 292466 77378 292702 77614
rect 292466 41698 292702 41934
rect 292466 41378 292702 41614
rect 292466 5698 292702 5934
rect 292466 5378 292702 5614
rect 292466 -2422 292702 -2186
rect 292466 -2742 292702 -2506
rect 295946 693178 296182 693414
rect 295946 692858 296182 693094
rect 295946 657178 296182 657414
rect 295946 656858 296182 657094
rect 295946 621178 296182 621414
rect 295946 620858 296182 621094
rect 295946 585178 296182 585414
rect 295946 584858 296182 585094
rect 295946 549178 296182 549414
rect 295946 548858 296182 549094
rect 295946 513178 296182 513414
rect 295946 512858 296182 513094
rect 295946 477178 296182 477414
rect 295946 476858 296182 477094
rect 295946 441178 296182 441414
rect 295946 440858 296182 441094
rect 295946 405178 296182 405414
rect 295946 404858 296182 405094
rect 295946 369178 296182 369414
rect 295946 368858 296182 369094
rect 295946 333178 296182 333414
rect 295946 332858 296182 333094
rect 295946 297178 296182 297414
rect 295946 296858 296182 297094
rect 295946 261178 296182 261414
rect 295946 260858 296182 261094
rect 295946 225178 296182 225414
rect 295946 224858 296182 225094
rect 295946 189178 296182 189414
rect 295946 188858 296182 189094
rect 295946 153178 296182 153414
rect 295946 152858 296182 153094
rect 295946 117178 296182 117414
rect 295946 116858 296182 117094
rect 295946 81178 296182 81414
rect 295946 80858 296182 81094
rect 295946 45178 296182 45414
rect 295946 44858 296182 45094
rect 295946 9178 296182 9414
rect 295946 8858 296182 9094
rect 295946 -4262 296182 -4026
rect 295946 -4582 296182 -4346
rect 317426 711042 317662 711278
rect 317426 710722 317662 710958
rect 313946 709202 314182 709438
rect 313946 708882 314182 709118
rect 310466 707362 310702 707598
rect 310466 707042 310702 707278
rect 299426 696658 299662 696894
rect 299426 696338 299662 696574
rect 299426 660658 299662 660894
rect 299426 660338 299662 660574
rect 299426 624658 299662 624894
rect 299426 624338 299662 624574
rect 299426 588658 299662 588894
rect 299426 588338 299662 588574
rect 299426 552658 299662 552894
rect 299426 552338 299662 552574
rect 299426 516658 299662 516894
rect 299426 516338 299662 516574
rect 299426 480658 299662 480894
rect 299426 480338 299662 480574
rect 299426 444658 299662 444894
rect 299426 444338 299662 444574
rect 299426 408658 299662 408894
rect 299426 408338 299662 408574
rect 299426 372658 299662 372894
rect 299426 372338 299662 372574
rect 299426 336658 299662 336894
rect 299426 336338 299662 336574
rect 299426 300658 299662 300894
rect 299426 300338 299662 300574
rect 299426 264658 299662 264894
rect 299426 264338 299662 264574
rect 299426 228658 299662 228894
rect 299426 228338 299662 228574
rect 299426 192658 299662 192894
rect 299426 192338 299662 192574
rect 299426 156658 299662 156894
rect 299426 156338 299662 156574
rect 299426 120658 299662 120894
rect 299426 120338 299662 120574
rect 299426 84658 299662 84894
rect 299426 84338 299662 84574
rect 299426 48658 299662 48894
rect 299426 48338 299662 48574
rect 299426 12658 299662 12894
rect 299426 12338 299662 12574
rect 281426 -7022 281662 -6786
rect 281426 -7342 281662 -7106
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310466 671698 310702 671934
rect 310466 671378 310702 671614
rect 310466 635698 310702 635934
rect 310466 635378 310702 635614
rect 310466 599698 310702 599934
rect 310466 599378 310702 599614
rect 310466 563698 310702 563934
rect 310466 563378 310702 563614
rect 310466 527698 310702 527934
rect 310466 527378 310702 527614
rect 310466 491698 310702 491934
rect 310466 491378 310702 491614
rect 310466 455698 310702 455934
rect 310466 455378 310702 455614
rect 310466 419698 310702 419934
rect 310466 419378 310702 419614
rect 310466 383698 310702 383934
rect 310466 383378 310702 383614
rect 310466 347698 310702 347934
rect 310466 347378 310702 347614
rect 310466 311698 310702 311934
rect 310466 311378 310702 311614
rect 310466 275698 310702 275934
rect 310466 275378 310702 275614
rect 310466 239698 310702 239934
rect 310466 239378 310702 239614
rect 310466 203698 310702 203934
rect 310466 203378 310702 203614
rect 310466 167698 310702 167934
rect 310466 167378 310702 167614
rect 310466 131698 310702 131934
rect 310466 131378 310702 131614
rect 310466 95698 310702 95934
rect 310466 95378 310702 95614
rect 310466 59698 310702 59934
rect 310466 59378 310702 59614
rect 310466 23698 310702 23934
rect 310466 23378 310702 23614
rect 310466 -3342 310702 -3106
rect 310466 -3662 310702 -3426
rect 313946 675178 314182 675414
rect 313946 674858 314182 675094
rect 313946 639178 314182 639414
rect 313946 638858 314182 639094
rect 313946 603178 314182 603414
rect 313946 602858 314182 603094
rect 313946 567178 314182 567414
rect 313946 566858 314182 567094
rect 313946 531178 314182 531414
rect 313946 530858 314182 531094
rect 313946 495178 314182 495414
rect 313946 494858 314182 495094
rect 313946 459178 314182 459414
rect 313946 458858 314182 459094
rect 313946 423178 314182 423414
rect 313946 422858 314182 423094
rect 313946 387178 314182 387414
rect 313946 386858 314182 387094
rect 313946 351178 314182 351414
rect 313946 350858 314182 351094
rect 313946 315178 314182 315414
rect 313946 314858 314182 315094
rect 313946 279178 314182 279414
rect 313946 278858 314182 279094
rect 313946 243178 314182 243414
rect 313946 242858 314182 243094
rect 313946 207178 314182 207414
rect 313946 206858 314182 207094
rect 313946 171178 314182 171414
rect 313946 170858 314182 171094
rect 313946 135178 314182 135414
rect 313946 134858 314182 135094
rect 313946 99178 314182 99414
rect 313946 98858 314182 99094
rect 313946 63178 314182 63414
rect 313946 62858 314182 63094
rect 313946 27178 314182 27414
rect 313946 26858 314182 27094
rect 313946 -5182 314182 -4946
rect 313946 -5502 314182 -5266
rect 335426 710122 335662 710358
rect 335426 709802 335662 710038
rect 331946 708282 332182 708518
rect 331946 707962 332182 708198
rect 328466 706442 328702 706678
rect 328466 706122 328702 706358
rect 317426 678658 317662 678894
rect 317426 678338 317662 678574
rect 317426 642658 317662 642894
rect 317426 642338 317662 642574
rect 317426 606658 317662 606894
rect 317426 606338 317662 606574
rect 317426 570658 317662 570894
rect 317426 570338 317662 570574
rect 317426 534658 317662 534894
rect 317426 534338 317662 534574
rect 317426 498658 317662 498894
rect 317426 498338 317662 498574
rect 317426 462658 317662 462894
rect 317426 462338 317662 462574
rect 317426 426658 317662 426894
rect 317426 426338 317662 426574
rect 317426 390658 317662 390894
rect 317426 390338 317662 390574
rect 317426 354658 317662 354894
rect 317426 354338 317662 354574
rect 317426 318658 317662 318894
rect 317426 318338 317662 318574
rect 317426 282658 317662 282894
rect 317426 282338 317662 282574
rect 317426 246658 317662 246894
rect 317426 246338 317662 246574
rect 317426 210658 317662 210894
rect 317426 210338 317662 210574
rect 317426 174658 317662 174894
rect 317426 174338 317662 174574
rect 317426 138658 317662 138894
rect 317426 138338 317662 138574
rect 317426 102658 317662 102894
rect 317426 102338 317662 102574
rect 317426 66658 317662 66894
rect 317426 66338 317662 66574
rect 317426 30658 317662 30894
rect 317426 30338 317662 30574
rect 299426 -6102 299662 -5866
rect 299426 -6422 299662 -6186
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328466 689698 328702 689934
rect 328466 689378 328702 689614
rect 328466 653698 328702 653934
rect 328466 653378 328702 653614
rect 328466 617698 328702 617934
rect 328466 617378 328702 617614
rect 328466 581698 328702 581934
rect 328466 581378 328702 581614
rect 328466 545698 328702 545934
rect 328466 545378 328702 545614
rect 328466 509698 328702 509934
rect 328466 509378 328702 509614
rect 328466 473698 328702 473934
rect 328466 473378 328702 473614
rect 328466 437698 328702 437934
rect 328466 437378 328702 437614
rect 328466 401698 328702 401934
rect 328466 401378 328702 401614
rect 328466 365698 328702 365934
rect 328466 365378 328702 365614
rect 328466 329698 328702 329934
rect 328466 329378 328702 329614
rect 328466 293698 328702 293934
rect 328466 293378 328702 293614
rect 328466 257698 328702 257934
rect 328466 257378 328702 257614
rect 328466 221698 328702 221934
rect 328466 221378 328702 221614
rect 328466 185698 328702 185934
rect 328466 185378 328702 185614
rect 328466 149698 328702 149934
rect 328466 149378 328702 149614
rect 328466 113698 328702 113934
rect 328466 113378 328702 113614
rect 328466 77698 328702 77934
rect 328466 77378 328702 77614
rect 328466 41698 328702 41934
rect 328466 41378 328702 41614
rect 328466 5698 328702 5934
rect 328466 5378 328702 5614
rect 328466 -2422 328702 -2186
rect 328466 -2742 328702 -2506
rect 331946 693178 332182 693414
rect 331946 692858 332182 693094
rect 331946 657178 332182 657414
rect 331946 656858 332182 657094
rect 331946 621178 332182 621414
rect 331946 620858 332182 621094
rect 331946 585178 332182 585414
rect 331946 584858 332182 585094
rect 331946 549178 332182 549414
rect 331946 548858 332182 549094
rect 331946 513178 332182 513414
rect 331946 512858 332182 513094
rect 331946 477178 332182 477414
rect 331946 476858 332182 477094
rect 331946 441178 332182 441414
rect 331946 440858 332182 441094
rect 331946 405178 332182 405414
rect 331946 404858 332182 405094
rect 331946 369178 332182 369414
rect 331946 368858 332182 369094
rect 331946 333178 332182 333414
rect 331946 332858 332182 333094
rect 331946 297178 332182 297414
rect 331946 296858 332182 297094
rect 331946 261178 332182 261414
rect 331946 260858 332182 261094
rect 331946 225178 332182 225414
rect 331946 224858 332182 225094
rect 331946 189178 332182 189414
rect 331946 188858 332182 189094
rect 331946 153178 332182 153414
rect 331946 152858 332182 153094
rect 331946 117178 332182 117414
rect 331946 116858 332182 117094
rect 331946 81178 332182 81414
rect 331946 80858 332182 81094
rect 331946 45178 332182 45414
rect 331946 44858 332182 45094
rect 331946 9178 332182 9414
rect 331946 8858 332182 9094
rect 331946 -4262 332182 -4026
rect 331946 -4582 332182 -4346
rect 353426 711042 353662 711278
rect 353426 710722 353662 710958
rect 349946 709202 350182 709438
rect 349946 708882 350182 709118
rect 346466 707362 346702 707598
rect 346466 707042 346702 707278
rect 335426 696658 335662 696894
rect 335426 696338 335662 696574
rect 335426 660658 335662 660894
rect 335426 660338 335662 660574
rect 335426 624658 335662 624894
rect 335426 624338 335662 624574
rect 335426 588658 335662 588894
rect 335426 588338 335662 588574
rect 335426 552658 335662 552894
rect 335426 552338 335662 552574
rect 335426 516658 335662 516894
rect 335426 516338 335662 516574
rect 335426 480658 335662 480894
rect 335426 480338 335662 480574
rect 335426 444658 335662 444894
rect 335426 444338 335662 444574
rect 335426 408658 335662 408894
rect 335426 408338 335662 408574
rect 335426 372658 335662 372894
rect 335426 372338 335662 372574
rect 335426 336658 335662 336894
rect 335426 336338 335662 336574
rect 335426 300658 335662 300894
rect 335426 300338 335662 300574
rect 335426 264658 335662 264894
rect 335426 264338 335662 264574
rect 335426 228658 335662 228894
rect 335426 228338 335662 228574
rect 335426 192658 335662 192894
rect 335426 192338 335662 192574
rect 335426 156658 335662 156894
rect 335426 156338 335662 156574
rect 335426 120658 335662 120894
rect 335426 120338 335662 120574
rect 335426 84658 335662 84894
rect 335426 84338 335662 84574
rect 335426 48658 335662 48894
rect 335426 48338 335662 48574
rect 335426 12658 335662 12894
rect 335426 12338 335662 12574
rect 317426 -7022 317662 -6786
rect 317426 -7342 317662 -7106
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 346466 671698 346702 671934
rect 346466 671378 346702 671614
rect 346466 635698 346702 635934
rect 346466 635378 346702 635614
rect 346466 599698 346702 599934
rect 346466 599378 346702 599614
rect 346466 563698 346702 563934
rect 346466 563378 346702 563614
rect 346466 527698 346702 527934
rect 346466 527378 346702 527614
rect 346466 491698 346702 491934
rect 346466 491378 346702 491614
rect 346466 455698 346702 455934
rect 346466 455378 346702 455614
rect 346466 419698 346702 419934
rect 346466 419378 346702 419614
rect 346466 383698 346702 383934
rect 346466 383378 346702 383614
rect 344790 363342 345026 363578
rect 344790 360622 345026 360858
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346466 347698 346702 347934
rect 346466 347378 346702 347614
rect 346466 311698 346702 311934
rect 346466 311378 346702 311614
rect 346466 275698 346702 275934
rect 346466 275378 346702 275614
rect 346466 239698 346702 239934
rect 346466 239378 346702 239614
rect 346466 203698 346702 203934
rect 346466 203378 346702 203614
rect 346466 167698 346702 167934
rect 346466 167378 346702 167614
rect 346466 131698 346702 131934
rect 346466 131378 346702 131614
rect 346466 95698 346702 95934
rect 346466 95378 346702 95614
rect 346466 59698 346702 59934
rect 346466 59378 346702 59614
rect 346466 23698 346702 23934
rect 346466 23378 346702 23614
rect 346466 -3342 346702 -3106
rect 346466 -3662 346702 -3426
rect 349946 675178 350182 675414
rect 349946 674858 350182 675094
rect 349946 639178 350182 639414
rect 349946 638858 350182 639094
rect 349946 603178 350182 603414
rect 349946 602858 350182 603094
rect 349946 567178 350182 567414
rect 349946 566858 350182 567094
rect 349946 531178 350182 531414
rect 349946 530858 350182 531094
rect 349946 495178 350182 495414
rect 349946 494858 350182 495094
rect 349946 459178 350182 459414
rect 349946 458858 350182 459094
rect 349946 423178 350182 423414
rect 349946 422858 350182 423094
rect 349946 387178 350182 387414
rect 349946 386858 350182 387094
rect 349946 351178 350182 351414
rect 349946 350858 350182 351094
rect 349946 315178 350182 315414
rect 349946 314858 350182 315094
rect 349946 279178 350182 279414
rect 349946 278858 350182 279094
rect 349946 243178 350182 243414
rect 349946 242858 350182 243094
rect 349946 207178 350182 207414
rect 349946 206858 350182 207094
rect 349946 171178 350182 171414
rect 349946 170858 350182 171094
rect 349946 135178 350182 135414
rect 349946 134858 350182 135094
rect 349946 99178 350182 99414
rect 349946 98858 350182 99094
rect 349946 63178 350182 63414
rect 349946 62858 350182 63094
rect 349946 27178 350182 27414
rect 349946 26858 350182 27094
rect 349946 -5182 350182 -4946
rect 349946 -5502 350182 -5266
rect 371426 710122 371662 710358
rect 371426 709802 371662 710038
rect 367946 708282 368182 708518
rect 367946 707962 368182 708198
rect 364466 706442 364702 706678
rect 364466 706122 364702 706358
rect 353426 678658 353662 678894
rect 353426 678338 353662 678574
rect 353426 642658 353662 642894
rect 353426 642338 353662 642574
rect 353426 606658 353662 606894
rect 353426 606338 353662 606574
rect 353426 570658 353662 570894
rect 353426 570338 353662 570574
rect 353426 534658 353662 534894
rect 353426 534338 353662 534574
rect 353426 498658 353662 498894
rect 353426 498338 353662 498574
rect 353426 462658 353662 462894
rect 353426 462338 353662 462574
rect 353426 426658 353662 426894
rect 353426 426338 353662 426574
rect 353426 390658 353662 390894
rect 353426 390338 353662 390574
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 359510 360622 359746 360858
rect 353426 354658 353662 354894
rect 353426 354338 353662 354574
rect 353426 318658 353662 318894
rect 353426 318338 353662 318574
rect 353426 282658 353662 282894
rect 353426 282338 353662 282574
rect 353426 246658 353662 246894
rect 353426 246338 353662 246574
rect 353426 210658 353662 210894
rect 353426 210338 353662 210574
rect 353426 174658 353662 174894
rect 353426 174338 353662 174574
rect 353426 138658 353662 138894
rect 353426 138338 353662 138574
rect 353426 102658 353662 102894
rect 353426 102338 353662 102574
rect 353426 66658 353662 66894
rect 353426 66338 353662 66574
rect 353426 30658 353662 30894
rect 353426 30338 353662 30574
rect 335426 -6102 335662 -5866
rect 335426 -6422 335662 -6186
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364466 689698 364702 689934
rect 364466 689378 364702 689614
rect 364466 653698 364702 653934
rect 364466 653378 364702 653614
rect 364466 617698 364702 617934
rect 364466 617378 364702 617614
rect 364466 581698 364702 581934
rect 364466 581378 364702 581614
rect 364466 545698 364702 545934
rect 364466 545378 364702 545614
rect 364466 509698 364702 509934
rect 364466 509378 364702 509614
rect 364466 473698 364702 473934
rect 364466 473378 364702 473614
rect 364466 437698 364702 437934
rect 364466 437378 364702 437614
rect 364466 401698 364702 401934
rect 364466 401378 364702 401614
rect 364466 365698 364702 365934
rect 364466 365378 364702 365614
rect 364466 329698 364702 329934
rect 364466 329378 364702 329614
rect 364466 293698 364702 293934
rect 364466 293378 364702 293614
rect 364466 257698 364702 257934
rect 364466 257378 364702 257614
rect 364466 221698 364702 221934
rect 364466 221378 364702 221614
rect 364466 185698 364702 185934
rect 364466 185378 364702 185614
rect 364466 149698 364702 149934
rect 364466 149378 364702 149614
rect 364466 113698 364702 113934
rect 364466 113378 364702 113614
rect 364466 77698 364702 77934
rect 364466 77378 364702 77614
rect 364466 41698 364702 41934
rect 364466 41378 364702 41614
rect 364466 5698 364702 5934
rect 364466 5378 364702 5614
rect 364466 -2422 364702 -2186
rect 364466 -2742 364702 -2506
rect 367946 693178 368182 693414
rect 367946 692858 368182 693094
rect 367946 657178 368182 657414
rect 367946 656858 368182 657094
rect 367946 621178 368182 621414
rect 367946 620858 368182 621094
rect 367946 585178 368182 585414
rect 367946 584858 368182 585094
rect 367946 549178 368182 549414
rect 367946 548858 368182 549094
rect 367946 513178 368182 513414
rect 367946 512858 368182 513094
rect 367946 477178 368182 477414
rect 367946 476858 368182 477094
rect 367946 441178 368182 441414
rect 367946 440858 368182 441094
rect 367946 405178 368182 405414
rect 367946 404858 368182 405094
rect 367946 369178 368182 369414
rect 367946 368858 368182 369094
rect 367946 333178 368182 333414
rect 367946 332858 368182 333094
rect 367946 297178 368182 297414
rect 367946 296858 368182 297094
rect 367946 261178 368182 261414
rect 367946 260858 368182 261094
rect 367946 225178 368182 225414
rect 367946 224858 368182 225094
rect 367946 189178 368182 189414
rect 367946 188858 368182 189094
rect 367946 153178 368182 153414
rect 367946 152858 368182 153094
rect 367946 117178 368182 117414
rect 367946 116858 368182 117094
rect 367946 81178 368182 81414
rect 367946 80858 368182 81094
rect 367946 45178 368182 45414
rect 367946 44858 368182 45094
rect 367946 9178 368182 9414
rect 367946 8858 368182 9094
rect 367946 -4262 368182 -4026
rect 367946 -4582 368182 -4346
rect 389426 711042 389662 711278
rect 389426 710722 389662 710958
rect 385946 709202 386182 709438
rect 385946 708882 386182 709118
rect 382466 707362 382702 707598
rect 382466 707042 382702 707278
rect 371426 696658 371662 696894
rect 371426 696338 371662 696574
rect 371426 660658 371662 660894
rect 371426 660338 371662 660574
rect 371426 624658 371662 624894
rect 371426 624338 371662 624574
rect 371426 588658 371662 588894
rect 371426 588338 371662 588574
rect 371426 552658 371662 552894
rect 371426 552338 371662 552574
rect 371426 516658 371662 516894
rect 371426 516338 371662 516574
rect 371426 480658 371662 480894
rect 371426 480338 371662 480574
rect 371426 444658 371662 444894
rect 371426 444338 371662 444574
rect 371426 408658 371662 408894
rect 371426 408338 371662 408574
rect 371426 372658 371662 372894
rect 371426 372338 371662 372574
rect 371426 336658 371662 336894
rect 371426 336338 371662 336574
rect 371426 300658 371662 300894
rect 371426 300338 371662 300574
rect 371426 264658 371662 264894
rect 371426 264338 371662 264574
rect 371426 228658 371662 228894
rect 371426 228338 371662 228574
rect 371426 192658 371662 192894
rect 371426 192338 371662 192574
rect 371426 156658 371662 156894
rect 371426 156338 371662 156574
rect 371426 120658 371662 120894
rect 371426 120338 371662 120574
rect 371426 84658 371662 84894
rect 371426 84338 371662 84574
rect 371426 48658 371662 48894
rect 371426 48338 371662 48574
rect 371426 12658 371662 12894
rect 371426 12338 371662 12574
rect 353426 -7022 353662 -6786
rect 353426 -7342 353662 -7106
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382466 671698 382702 671934
rect 382466 671378 382702 671614
rect 382466 635698 382702 635934
rect 382466 635378 382702 635614
rect 382466 599698 382702 599934
rect 382466 599378 382702 599614
rect 382466 563698 382702 563934
rect 382466 563378 382702 563614
rect 382466 527698 382702 527934
rect 382466 527378 382702 527614
rect 382466 491698 382702 491934
rect 382466 491378 382702 491614
rect 382466 455698 382702 455934
rect 382466 455378 382702 455614
rect 382466 419698 382702 419934
rect 382466 419378 382702 419614
rect 382466 383698 382702 383934
rect 382466 383378 382702 383614
rect 382466 347698 382702 347934
rect 382466 347378 382702 347614
rect 382466 311698 382702 311934
rect 382466 311378 382702 311614
rect 382466 275698 382702 275934
rect 382466 275378 382702 275614
rect 382466 239698 382702 239934
rect 382466 239378 382702 239614
rect 382466 203698 382702 203934
rect 382466 203378 382702 203614
rect 382466 167698 382702 167934
rect 382466 167378 382702 167614
rect 382466 131698 382702 131934
rect 382466 131378 382702 131614
rect 382466 95698 382702 95934
rect 382466 95378 382702 95614
rect 382466 59698 382702 59934
rect 382466 59378 382702 59614
rect 382466 23698 382702 23934
rect 382466 23378 382702 23614
rect 382466 -3342 382702 -3106
rect 382466 -3662 382702 -3426
rect 385946 675178 386182 675414
rect 385946 674858 386182 675094
rect 385946 639178 386182 639414
rect 385946 638858 386182 639094
rect 385946 603178 386182 603414
rect 385946 602858 386182 603094
rect 385946 567178 386182 567414
rect 385946 566858 386182 567094
rect 385946 531178 386182 531414
rect 385946 530858 386182 531094
rect 385946 495178 386182 495414
rect 385946 494858 386182 495094
rect 385946 459178 386182 459414
rect 385946 458858 386182 459094
rect 385946 423178 386182 423414
rect 385946 422858 386182 423094
rect 385946 387178 386182 387414
rect 385946 386858 386182 387094
rect 385946 351178 386182 351414
rect 385946 350858 386182 351094
rect 385946 315178 386182 315414
rect 385946 314858 386182 315094
rect 385946 279178 386182 279414
rect 385946 278858 386182 279094
rect 385946 243178 386182 243414
rect 385946 242858 386182 243094
rect 385946 207178 386182 207414
rect 385946 206858 386182 207094
rect 385946 171178 386182 171414
rect 385946 170858 386182 171094
rect 385946 135178 386182 135414
rect 385946 134858 386182 135094
rect 385946 99178 386182 99414
rect 385946 98858 386182 99094
rect 385946 63178 386182 63414
rect 385946 62858 386182 63094
rect 385946 27178 386182 27414
rect 385946 26858 386182 27094
rect 385946 -5182 386182 -4946
rect 385946 -5502 386182 -5266
rect 407426 710122 407662 710358
rect 407426 709802 407662 710038
rect 403946 708282 404182 708518
rect 403946 707962 404182 708198
rect 400466 706442 400702 706678
rect 400466 706122 400702 706358
rect 389426 678658 389662 678894
rect 389426 678338 389662 678574
rect 389426 642658 389662 642894
rect 389426 642338 389662 642574
rect 389426 606658 389662 606894
rect 389426 606338 389662 606574
rect 389426 570658 389662 570894
rect 389426 570338 389662 570574
rect 389426 534658 389662 534894
rect 389426 534338 389662 534574
rect 389426 498658 389662 498894
rect 389426 498338 389662 498574
rect 389426 462658 389662 462894
rect 389426 462338 389662 462574
rect 389426 426658 389662 426894
rect 389426 426338 389662 426574
rect 389426 390658 389662 390894
rect 389426 390338 389662 390574
rect 389426 354658 389662 354894
rect 389426 354338 389662 354574
rect 389426 318658 389662 318894
rect 389426 318338 389662 318574
rect 389426 282658 389662 282894
rect 389426 282338 389662 282574
rect 389426 246658 389662 246894
rect 389426 246338 389662 246574
rect 389426 210658 389662 210894
rect 389426 210338 389662 210574
rect 389426 174658 389662 174894
rect 389426 174338 389662 174574
rect 389426 138658 389662 138894
rect 389426 138338 389662 138574
rect 389426 102658 389662 102894
rect 389426 102338 389662 102574
rect 389426 66658 389662 66894
rect 389426 66338 389662 66574
rect 389426 30658 389662 30894
rect 389426 30338 389662 30574
rect 371426 -6102 371662 -5866
rect 371426 -6422 371662 -6186
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400466 689698 400702 689934
rect 400466 689378 400702 689614
rect 400466 653698 400702 653934
rect 400466 653378 400702 653614
rect 400466 617698 400702 617934
rect 400466 617378 400702 617614
rect 400466 581698 400702 581934
rect 400466 581378 400702 581614
rect 400466 545698 400702 545934
rect 400466 545378 400702 545614
rect 400466 509698 400702 509934
rect 400466 509378 400702 509614
rect 400466 473698 400702 473934
rect 400466 473378 400702 473614
rect 400466 437698 400702 437934
rect 400466 437378 400702 437614
rect 400466 401698 400702 401934
rect 400466 401378 400702 401614
rect 400466 365698 400702 365934
rect 400466 365378 400702 365614
rect 400466 329698 400702 329934
rect 400466 329378 400702 329614
rect 400466 293698 400702 293934
rect 400466 293378 400702 293614
rect 400466 257698 400702 257934
rect 400466 257378 400702 257614
rect 400466 221698 400702 221934
rect 400466 221378 400702 221614
rect 400466 185698 400702 185934
rect 400466 185378 400702 185614
rect 400466 149698 400702 149934
rect 400466 149378 400702 149614
rect 400466 113698 400702 113934
rect 400466 113378 400702 113614
rect 400466 77698 400702 77934
rect 400466 77378 400702 77614
rect 400466 41698 400702 41934
rect 400466 41378 400702 41614
rect 400466 5698 400702 5934
rect 400466 5378 400702 5614
rect 400466 -2422 400702 -2186
rect 400466 -2742 400702 -2506
rect 403946 693178 404182 693414
rect 403946 692858 404182 693094
rect 403946 657178 404182 657414
rect 403946 656858 404182 657094
rect 403946 621178 404182 621414
rect 403946 620858 404182 621094
rect 403946 585178 404182 585414
rect 403946 584858 404182 585094
rect 403946 549178 404182 549414
rect 403946 548858 404182 549094
rect 403946 513178 404182 513414
rect 403946 512858 404182 513094
rect 403946 477178 404182 477414
rect 403946 476858 404182 477094
rect 403946 441178 404182 441414
rect 403946 440858 404182 441094
rect 403946 405178 404182 405414
rect 403946 404858 404182 405094
rect 403946 369178 404182 369414
rect 403946 368858 404182 369094
rect 403946 333178 404182 333414
rect 403946 332858 404182 333094
rect 403946 297178 404182 297414
rect 403946 296858 404182 297094
rect 403946 261178 404182 261414
rect 403946 260858 404182 261094
rect 403946 225178 404182 225414
rect 403946 224858 404182 225094
rect 403946 189178 404182 189414
rect 403946 188858 404182 189094
rect 403946 153178 404182 153414
rect 403946 152858 404182 153094
rect 403946 117178 404182 117414
rect 403946 116858 404182 117094
rect 403946 81178 404182 81414
rect 403946 80858 404182 81094
rect 403946 45178 404182 45414
rect 403946 44858 404182 45094
rect 403946 9178 404182 9414
rect 403946 8858 404182 9094
rect 403946 -4262 404182 -4026
rect 403946 -4582 404182 -4346
rect 425426 711042 425662 711278
rect 425426 710722 425662 710958
rect 421946 709202 422182 709438
rect 421946 708882 422182 709118
rect 418466 707362 418702 707598
rect 418466 707042 418702 707278
rect 407426 696658 407662 696894
rect 407426 696338 407662 696574
rect 407426 660658 407662 660894
rect 407426 660338 407662 660574
rect 407426 624658 407662 624894
rect 407426 624338 407662 624574
rect 407426 588658 407662 588894
rect 407426 588338 407662 588574
rect 407426 552658 407662 552894
rect 407426 552338 407662 552574
rect 407426 516658 407662 516894
rect 407426 516338 407662 516574
rect 407426 480658 407662 480894
rect 407426 480338 407662 480574
rect 407426 444658 407662 444894
rect 407426 444338 407662 444574
rect 407426 408658 407662 408894
rect 407426 408338 407662 408574
rect 407426 372658 407662 372894
rect 407426 372338 407662 372574
rect 407426 336658 407662 336894
rect 407426 336338 407662 336574
rect 407426 300658 407662 300894
rect 407426 300338 407662 300574
rect 407426 264658 407662 264894
rect 407426 264338 407662 264574
rect 407426 228658 407662 228894
rect 407426 228338 407662 228574
rect 407426 192658 407662 192894
rect 407426 192338 407662 192574
rect 407426 156658 407662 156894
rect 407426 156338 407662 156574
rect 407426 120658 407662 120894
rect 407426 120338 407662 120574
rect 407426 84658 407662 84894
rect 407426 84338 407662 84574
rect 407426 48658 407662 48894
rect 407426 48338 407662 48574
rect 407426 12658 407662 12894
rect 407426 12338 407662 12574
rect 389426 -7022 389662 -6786
rect 389426 -7342 389662 -7106
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418466 671698 418702 671934
rect 418466 671378 418702 671614
rect 418466 635698 418702 635934
rect 418466 635378 418702 635614
rect 418466 599698 418702 599934
rect 418466 599378 418702 599614
rect 418466 563698 418702 563934
rect 418466 563378 418702 563614
rect 418466 527698 418702 527934
rect 418466 527378 418702 527614
rect 418466 491698 418702 491934
rect 418466 491378 418702 491614
rect 418466 455698 418702 455934
rect 418466 455378 418702 455614
rect 418466 419698 418702 419934
rect 418466 419378 418702 419614
rect 418466 383698 418702 383934
rect 418466 383378 418702 383614
rect 418466 347698 418702 347934
rect 418466 347378 418702 347614
rect 418466 311698 418702 311934
rect 418466 311378 418702 311614
rect 418466 275698 418702 275934
rect 418466 275378 418702 275614
rect 418466 239698 418702 239934
rect 418466 239378 418702 239614
rect 418466 203698 418702 203934
rect 418466 203378 418702 203614
rect 418466 167698 418702 167934
rect 418466 167378 418702 167614
rect 418466 131698 418702 131934
rect 418466 131378 418702 131614
rect 418466 95698 418702 95934
rect 418466 95378 418702 95614
rect 418466 59698 418702 59934
rect 418466 59378 418702 59614
rect 418466 23698 418702 23934
rect 418466 23378 418702 23614
rect 418466 -3342 418702 -3106
rect 418466 -3662 418702 -3426
rect 421946 675178 422182 675414
rect 421946 674858 422182 675094
rect 421946 639178 422182 639414
rect 421946 638858 422182 639094
rect 421946 603178 422182 603414
rect 421946 602858 422182 603094
rect 421946 567178 422182 567414
rect 421946 566858 422182 567094
rect 421946 531178 422182 531414
rect 421946 530858 422182 531094
rect 421946 495178 422182 495414
rect 421946 494858 422182 495094
rect 421946 459178 422182 459414
rect 421946 458858 422182 459094
rect 421946 423178 422182 423414
rect 421946 422858 422182 423094
rect 421946 387178 422182 387414
rect 421946 386858 422182 387094
rect 421946 351178 422182 351414
rect 421946 350858 422182 351094
rect 421946 315178 422182 315414
rect 421946 314858 422182 315094
rect 421946 279178 422182 279414
rect 421946 278858 422182 279094
rect 421946 243178 422182 243414
rect 421946 242858 422182 243094
rect 421946 207178 422182 207414
rect 421946 206858 422182 207094
rect 421946 171178 422182 171414
rect 421946 170858 422182 171094
rect 421946 135178 422182 135414
rect 421946 134858 422182 135094
rect 421946 99178 422182 99414
rect 421946 98858 422182 99094
rect 421946 63178 422182 63414
rect 421946 62858 422182 63094
rect 421946 27178 422182 27414
rect 421946 26858 422182 27094
rect 421946 -5182 422182 -4946
rect 421946 -5502 422182 -5266
rect 443426 710122 443662 710358
rect 443426 709802 443662 710038
rect 439946 708282 440182 708518
rect 439946 707962 440182 708198
rect 436466 706442 436702 706678
rect 436466 706122 436702 706358
rect 425426 678658 425662 678894
rect 425426 678338 425662 678574
rect 425426 642658 425662 642894
rect 425426 642338 425662 642574
rect 425426 606658 425662 606894
rect 425426 606338 425662 606574
rect 425426 570658 425662 570894
rect 425426 570338 425662 570574
rect 425426 534658 425662 534894
rect 425426 534338 425662 534574
rect 425426 498658 425662 498894
rect 425426 498338 425662 498574
rect 425426 462658 425662 462894
rect 425426 462338 425662 462574
rect 425426 426658 425662 426894
rect 425426 426338 425662 426574
rect 425426 390658 425662 390894
rect 425426 390338 425662 390574
rect 425426 354658 425662 354894
rect 425426 354338 425662 354574
rect 425426 318658 425662 318894
rect 425426 318338 425662 318574
rect 425426 282658 425662 282894
rect 425426 282338 425662 282574
rect 425426 246658 425662 246894
rect 425426 246338 425662 246574
rect 425426 210658 425662 210894
rect 425426 210338 425662 210574
rect 425426 174658 425662 174894
rect 425426 174338 425662 174574
rect 425426 138658 425662 138894
rect 425426 138338 425662 138574
rect 425426 102658 425662 102894
rect 425426 102338 425662 102574
rect 425426 66658 425662 66894
rect 425426 66338 425662 66574
rect 425426 30658 425662 30894
rect 425426 30338 425662 30574
rect 407426 -6102 407662 -5866
rect 407426 -6422 407662 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436466 689698 436702 689934
rect 436466 689378 436702 689614
rect 436466 653698 436702 653934
rect 436466 653378 436702 653614
rect 436466 617698 436702 617934
rect 436466 617378 436702 617614
rect 436466 581698 436702 581934
rect 436466 581378 436702 581614
rect 436466 545698 436702 545934
rect 436466 545378 436702 545614
rect 436466 509698 436702 509934
rect 436466 509378 436702 509614
rect 436466 473698 436702 473934
rect 436466 473378 436702 473614
rect 436466 437698 436702 437934
rect 436466 437378 436702 437614
rect 436466 401698 436702 401934
rect 436466 401378 436702 401614
rect 436466 365698 436702 365934
rect 436466 365378 436702 365614
rect 436466 329698 436702 329934
rect 436466 329378 436702 329614
rect 436466 293698 436702 293934
rect 436466 293378 436702 293614
rect 436466 257698 436702 257934
rect 436466 257378 436702 257614
rect 436466 221698 436702 221934
rect 436466 221378 436702 221614
rect 436466 185698 436702 185934
rect 436466 185378 436702 185614
rect 436466 149698 436702 149934
rect 436466 149378 436702 149614
rect 436466 113698 436702 113934
rect 436466 113378 436702 113614
rect 436466 77698 436702 77934
rect 436466 77378 436702 77614
rect 436466 41698 436702 41934
rect 436466 41378 436702 41614
rect 436466 5698 436702 5934
rect 436466 5378 436702 5614
rect 436466 -2422 436702 -2186
rect 436466 -2742 436702 -2506
rect 439946 693178 440182 693414
rect 439946 692858 440182 693094
rect 439946 657178 440182 657414
rect 439946 656858 440182 657094
rect 439946 621178 440182 621414
rect 439946 620858 440182 621094
rect 439946 585178 440182 585414
rect 439946 584858 440182 585094
rect 439946 549178 440182 549414
rect 439946 548858 440182 549094
rect 439946 513178 440182 513414
rect 439946 512858 440182 513094
rect 439946 477178 440182 477414
rect 439946 476858 440182 477094
rect 439946 441178 440182 441414
rect 439946 440858 440182 441094
rect 439946 405178 440182 405414
rect 439946 404858 440182 405094
rect 439946 369178 440182 369414
rect 439946 368858 440182 369094
rect 439946 333178 440182 333414
rect 439946 332858 440182 333094
rect 439946 297178 440182 297414
rect 439946 296858 440182 297094
rect 439946 261178 440182 261414
rect 439946 260858 440182 261094
rect 439946 225178 440182 225414
rect 439946 224858 440182 225094
rect 439946 189178 440182 189414
rect 439946 188858 440182 189094
rect 439946 153178 440182 153414
rect 439946 152858 440182 153094
rect 439946 117178 440182 117414
rect 439946 116858 440182 117094
rect 439946 81178 440182 81414
rect 439946 80858 440182 81094
rect 439946 45178 440182 45414
rect 439946 44858 440182 45094
rect 439946 9178 440182 9414
rect 439946 8858 440182 9094
rect 439946 -4262 440182 -4026
rect 439946 -4582 440182 -4346
rect 461426 711042 461662 711278
rect 461426 710722 461662 710958
rect 457946 709202 458182 709438
rect 457946 708882 458182 709118
rect 454466 707362 454702 707598
rect 454466 707042 454702 707278
rect 443426 696658 443662 696894
rect 443426 696338 443662 696574
rect 443426 660658 443662 660894
rect 443426 660338 443662 660574
rect 443426 624658 443662 624894
rect 443426 624338 443662 624574
rect 443426 588658 443662 588894
rect 443426 588338 443662 588574
rect 443426 552658 443662 552894
rect 443426 552338 443662 552574
rect 443426 516658 443662 516894
rect 443426 516338 443662 516574
rect 443426 480658 443662 480894
rect 443426 480338 443662 480574
rect 443426 444658 443662 444894
rect 443426 444338 443662 444574
rect 443426 408658 443662 408894
rect 443426 408338 443662 408574
rect 443426 372658 443662 372894
rect 443426 372338 443662 372574
rect 443426 336658 443662 336894
rect 443426 336338 443662 336574
rect 443426 300658 443662 300894
rect 443426 300338 443662 300574
rect 443426 264658 443662 264894
rect 443426 264338 443662 264574
rect 443426 228658 443662 228894
rect 443426 228338 443662 228574
rect 443426 192658 443662 192894
rect 443426 192338 443662 192574
rect 443426 156658 443662 156894
rect 443426 156338 443662 156574
rect 443426 120658 443662 120894
rect 443426 120338 443662 120574
rect 443426 84658 443662 84894
rect 443426 84338 443662 84574
rect 443426 48658 443662 48894
rect 443426 48338 443662 48574
rect 443426 12658 443662 12894
rect 443426 12338 443662 12574
rect 425426 -7022 425662 -6786
rect 425426 -7342 425662 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454466 671698 454702 671934
rect 454466 671378 454702 671614
rect 454466 635698 454702 635934
rect 454466 635378 454702 635614
rect 454466 599698 454702 599934
rect 454466 599378 454702 599614
rect 454466 563698 454702 563934
rect 454466 563378 454702 563614
rect 454466 527698 454702 527934
rect 454466 527378 454702 527614
rect 454466 491698 454702 491934
rect 454466 491378 454702 491614
rect 454466 455698 454702 455934
rect 454466 455378 454702 455614
rect 454466 419698 454702 419934
rect 454466 419378 454702 419614
rect 454466 383698 454702 383934
rect 454466 383378 454702 383614
rect 454466 347698 454702 347934
rect 454466 347378 454702 347614
rect 454466 311698 454702 311934
rect 454466 311378 454702 311614
rect 454466 275698 454702 275934
rect 454466 275378 454702 275614
rect 454466 239698 454702 239934
rect 454466 239378 454702 239614
rect 454466 203698 454702 203934
rect 454466 203378 454702 203614
rect 454466 167698 454702 167934
rect 454466 167378 454702 167614
rect 454466 131698 454702 131934
rect 454466 131378 454702 131614
rect 454466 95698 454702 95934
rect 454466 95378 454702 95614
rect 454466 59698 454702 59934
rect 454466 59378 454702 59614
rect 454466 23698 454702 23934
rect 454466 23378 454702 23614
rect 454466 -3342 454702 -3106
rect 454466 -3662 454702 -3426
rect 457946 675178 458182 675414
rect 457946 674858 458182 675094
rect 457946 639178 458182 639414
rect 457946 638858 458182 639094
rect 457946 603178 458182 603414
rect 457946 602858 458182 603094
rect 457946 567178 458182 567414
rect 457946 566858 458182 567094
rect 457946 531178 458182 531414
rect 457946 530858 458182 531094
rect 457946 495178 458182 495414
rect 457946 494858 458182 495094
rect 457946 459178 458182 459414
rect 457946 458858 458182 459094
rect 457946 423178 458182 423414
rect 457946 422858 458182 423094
rect 457946 387178 458182 387414
rect 457946 386858 458182 387094
rect 457946 351178 458182 351414
rect 457946 350858 458182 351094
rect 457946 315178 458182 315414
rect 457946 314858 458182 315094
rect 457946 279178 458182 279414
rect 457946 278858 458182 279094
rect 457946 243178 458182 243414
rect 457946 242858 458182 243094
rect 457946 207178 458182 207414
rect 457946 206858 458182 207094
rect 457946 171178 458182 171414
rect 457946 170858 458182 171094
rect 457946 135178 458182 135414
rect 457946 134858 458182 135094
rect 457946 99178 458182 99414
rect 457946 98858 458182 99094
rect 457946 63178 458182 63414
rect 457946 62858 458182 63094
rect 457946 27178 458182 27414
rect 457946 26858 458182 27094
rect 457946 -5182 458182 -4946
rect 457946 -5502 458182 -5266
rect 479426 710122 479662 710358
rect 479426 709802 479662 710038
rect 475946 708282 476182 708518
rect 475946 707962 476182 708198
rect 472466 706442 472702 706678
rect 472466 706122 472702 706358
rect 461426 678658 461662 678894
rect 461426 678338 461662 678574
rect 461426 642658 461662 642894
rect 461426 642338 461662 642574
rect 461426 606658 461662 606894
rect 461426 606338 461662 606574
rect 461426 570658 461662 570894
rect 461426 570338 461662 570574
rect 461426 534658 461662 534894
rect 461426 534338 461662 534574
rect 461426 498658 461662 498894
rect 461426 498338 461662 498574
rect 461426 462658 461662 462894
rect 461426 462338 461662 462574
rect 461426 426658 461662 426894
rect 461426 426338 461662 426574
rect 461426 390658 461662 390894
rect 461426 390338 461662 390574
rect 461426 354658 461662 354894
rect 461426 354338 461662 354574
rect 461426 318658 461662 318894
rect 461426 318338 461662 318574
rect 461426 282658 461662 282894
rect 461426 282338 461662 282574
rect 461426 246658 461662 246894
rect 461426 246338 461662 246574
rect 461426 210658 461662 210894
rect 461426 210338 461662 210574
rect 461426 174658 461662 174894
rect 461426 174338 461662 174574
rect 461426 138658 461662 138894
rect 461426 138338 461662 138574
rect 461426 102658 461662 102894
rect 461426 102338 461662 102574
rect 461426 66658 461662 66894
rect 461426 66338 461662 66574
rect 461426 30658 461662 30894
rect 461426 30338 461662 30574
rect 443426 -6102 443662 -5866
rect 443426 -6422 443662 -6186
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472466 689698 472702 689934
rect 472466 689378 472702 689614
rect 472466 653698 472702 653934
rect 472466 653378 472702 653614
rect 472466 617698 472702 617934
rect 472466 617378 472702 617614
rect 472466 581698 472702 581934
rect 472466 581378 472702 581614
rect 472466 545698 472702 545934
rect 472466 545378 472702 545614
rect 472466 509698 472702 509934
rect 472466 509378 472702 509614
rect 472466 473698 472702 473934
rect 472466 473378 472702 473614
rect 472466 437698 472702 437934
rect 472466 437378 472702 437614
rect 472466 401698 472702 401934
rect 472466 401378 472702 401614
rect 472466 365698 472702 365934
rect 472466 365378 472702 365614
rect 472466 329698 472702 329934
rect 472466 329378 472702 329614
rect 472466 293698 472702 293934
rect 472466 293378 472702 293614
rect 472466 257698 472702 257934
rect 472466 257378 472702 257614
rect 472466 221698 472702 221934
rect 472466 221378 472702 221614
rect 472466 185698 472702 185934
rect 472466 185378 472702 185614
rect 472466 149698 472702 149934
rect 472466 149378 472702 149614
rect 472466 113698 472702 113934
rect 472466 113378 472702 113614
rect 472466 77698 472702 77934
rect 472466 77378 472702 77614
rect 472466 41698 472702 41934
rect 472466 41378 472702 41614
rect 472466 5698 472702 5934
rect 472466 5378 472702 5614
rect 472466 -2422 472702 -2186
rect 472466 -2742 472702 -2506
rect 475946 693178 476182 693414
rect 475946 692858 476182 693094
rect 475946 657178 476182 657414
rect 475946 656858 476182 657094
rect 475946 621178 476182 621414
rect 475946 620858 476182 621094
rect 475946 585178 476182 585414
rect 475946 584858 476182 585094
rect 475946 549178 476182 549414
rect 475946 548858 476182 549094
rect 475946 513178 476182 513414
rect 475946 512858 476182 513094
rect 475946 477178 476182 477414
rect 475946 476858 476182 477094
rect 475946 441178 476182 441414
rect 475946 440858 476182 441094
rect 475946 405178 476182 405414
rect 475946 404858 476182 405094
rect 475946 369178 476182 369414
rect 475946 368858 476182 369094
rect 475946 333178 476182 333414
rect 475946 332858 476182 333094
rect 475946 297178 476182 297414
rect 475946 296858 476182 297094
rect 475946 261178 476182 261414
rect 475946 260858 476182 261094
rect 475946 225178 476182 225414
rect 475946 224858 476182 225094
rect 475946 189178 476182 189414
rect 475946 188858 476182 189094
rect 475946 153178 476182 153414
rect 475946 152858 476182 153094
rect 475946 117178 476182 117414
rect 475946 116858 476182 117094
rect 475946 81178 476182 81414
rect 475946 80858 476182 81094
rect 475946 45178 476182 45414
rect 475946 44858 476182 45094
rect 475946 9178 476182 9414
rect 475946 8858 476182 9094
rect 475946 -4262 476182 -4026
rect 475946 -4582 476182 -4346
rect 497426 711042 497662 711278
rect 497426 710722 497662 710958
rect 493946 709202 494182 709438
rect 493946 708882 494182 709118
rect 490466 707362 490702 707598
rect 490466 707042 490702 707278
rect 479426 696658 479662 696894
rect 479426 696338 479662 696574
rect 479426 660658 479662 660894
rect 479426 660338 479662 660574
rect 479426 624658 479662 624894
rect 479426 624338 479662 624574
rect 479426 588658 479662 588894
rect 479426 588338 479662 588574
rect 479426 552658 479662 552894
rect 479426 552338 479662 552574
rect 479426 516658 479662 516894
rect 479426 516338 479662 516574
rect 479426 480658 479662 480894
rect 479426 480338 479662 480574
rect 479426 444658 479662 444894
rect 479426 444338 479662 444574
rect 479426 408658 479662 408894
rect 479426 408338 479662 408574
rect 479426 372658 479662 372894
rect 479426 372338 479662 372574
rect 479426 336658 479662 336894
rect 479426 336338 479662 336574
rect 479426 300658 479662 300894
rect 479426 300338 479662 300574
rect 479426 264658 479662 264894
rect 479426 264338 479662 264574
rect 479426 228658 479662 228894
rect 479426 228338 479662 228574
rect 479426 192658 479662 192894
rect 479426 192338 479662 192574
rect 479426 156658 479662 156894
rect 479426 156338 479662 156574
rect 479426 120658 479662 120894
rect 479426 120338 479662 120574
rect 479426 84658 479662 84894
rect 479426 84338 479662 84574
rect 479426 48658 479662 48894
rect 479426 48338 479662 48574
rect 479426 12658 479662 12894
rect 479426 12338 479662 12574
rect 461426 -7022 461662 -6786
rect 461426 -7342 461662 -7106
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490466 671698 490702 671934
rect 490466 671378 490702 671614
rect 490466 635698 490702 635934
rect 490466 635378 490702 635614
rect 490466 599698 490702 599934
rect 490466 599378 490702 599614
rect 490466 563698 490702 563934
rect 490466 563378 490702 563614
rect 490466 527698 490702 527934
rect 490466 527378 490702 527614
rect 490466 491698 490702 491934
rect 490466 491378 490702 491614
rect 490466 455698 490702 455934
rect 490466 455378 490702 455614
rect 490466 419698 490702 419934
rect 490466 419378 490702 419614
rect 490466 383698 490702 383934
rect 490466 383378 490702 383614
rect 490466 347698 490702 347934
rect 490466 347378 490702 347614
rect 490466 311698 490702 311934
rect 490466 311378 490702 311614
rect 490466 275698 490702 275934
rect 490466 275378 490702 275614
rect 490466 239698 490702 239934
rect 490466 239378 490702 239614
rect 490466 203698 490702 203934
rect 490466 203378 490702 203614
rect 490466 167698 490702 167934
rect 490466 167378 490702 167614
rect 490466 131698 490702 131934
rect 490466 131378 490702 131614
rect 490466 95698 490702 95934
rect 490466 95378 490702 95614
rect 490466 59698 490702 59934
rect 490466 59378 490702 59614
rect 490466 23698 490702 23934
rect 490466 23378 490702 23614
rect 490466 -3342 490702 -3106
rect 490466 -3662 490702 -3426
rect 493946 675178 494182 675414
rect 493946 674858 494182 675094
rect 493946 639178 494182 639414
rect 493946 638858 494182 639094
rect 493946 603178 494182 603414
rect 493946 602858 494182 603094
rect 493946 567178 494182 567414
rect 493946 566858 494182 567094
rect 493946 531178 494182 531414
rect 493946 530858 494182 531094
rect 493946 495178 494182 495414
rect 493946 494858 494182 495094
rect 493946 459178 494182 459414
rect 493946 458858 494182 459094
rect 493946 423178 494182 423414
rect 493946 422858 494182 423094
rect 493946 387178 494182 387414
rect 493946 386858 494182 387094
rect 493946 351178 494182 351414
rect 493946 350858 494182 351094
rect 493946 315178 494182 315414
rect 493946 314858 494182 315094
rect 493946 279178 494182 279414
rect 493946 278858 494182 279094
rect 493946 243178 494182 243414
rect 493946 242858 494182 243094
rect 493946 207178 494182 207414
rect 493946 206858 494182 207094
rect 493946 171178 494182 171414
rect 493946 170858 494182 171094
rect 493946 135178 494182 135414
rect 493946 134858 494182 135094
rect 493946 99178 494182 99414
rect 493946 98858 494182 99094
rect 493946 63178 494182 63414
rect 493946 62858 494182 63094
rect 493946 27178 494182 27414
rect 493946 26858 494182 27094
rect 493946 -5182 494182 -4946
rect 493946 -5502 494182 -5266
rect 515426 710122 515662 710358
rect 515426 709802 515662 710038
rect 511946 708282 512182 708518
rect 511946 707962 512182 708198
rect 508466 706442 508702 706678
rect 508466 706122 508702 706358
rect 497426 678658 497662 678894
rect 497426 678338 497662 678574
rect 497426 642658 497662 642894
rect 497426 642338 497662 642574
rect 497426 606658 497662 606894
rect 497426 606338 497662 606574
rect 497426 570658 497662 570894
rect 497426 570338 497662 570574
rect 497426 534658 497662 534894
rect 497426 534338 497662 534574
rect 497426 498658 497662 498894
rect 497426 498338 497662 498574
rect 497426 462658 497662 462894
rect 497426 462338 497662 462574
rect 497426 426658 497662 426894
rect 497426 426338 497662 426574
rect 497426 390658 497662 390894
rect 497426 390338 497662 390574
rect 497426 354658 497662 354894
rect 497426 354338 497662 354574
rect 497426 318658 497662 318894
rect 497426 318338 497662 318574
rect 497426 282658 497662 282894
rect 497426 282338 497662 282574
rect 497426 246658 497662 246894
rect 497426 246338 497662 246574
rect 497426 210658 497662 210894
rect 497426 210338 497662 210574
rect 497426 174658 497662 174894
rect 497426 174338 497662 174574
rect 497426 138658 497662 138894
rect 497426 138338 497662 138574
rect 497426 102658 497662 102894
rect 497426 102338 497662 102574
rect 497426 66658 497662 66894
rect 497426 66338 497662 66574
rect 497426 30658 497662 30894
rect 497426 30338 497662 30574
rect 479426 -6102 479662 -5866
rect 479426 -6422 479662 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508466 689698 508702 689934
rect 508466 689378 508702 689614
rect 508466 653698 508702 653934
rect 508466 653378 508702 653614
rect 508466 617698 508702 617934
rect 508466 617378 508702 617614
rect 508466 581698 508702 581934
rect 508466 581378 508702 581614
rect 508466 545698 508702 545934
rect 508466 545378 508702 545614
rect 508466 509698 508702 509934
rect 508466 509378 508702 509614
rect 508466 473698 508702 473934
rect 508466 473378 508702 473614
rect 508466 437698 508702 437934
rect 508466 437378 508702 437614
rect 508466 401698 508702 401934
rect 508466 401378 508702 401614
rect 508466 365698 508702 365934
rect 508466 365378 508702 365614
rect 508466 329698 508702 329934
rect 508466 329378 508702 329614
rect 508466 293698 508702 293934
rect 508466 293378 508702 293614
rect 508466 257698 508702 257934
rect 508466 257378 508702 257614
rect 508466 221698 508702 221934
rect 508466 221378 508702 221614
rect 508466 185698 508702 185934
rect 508466 185378 508702 185614
rect 508466 149698 508702 149934
rect 508466 149378 508702 149614
rect 508466 113698 508702 113934
rect 508466 113378 508702 113614
rect 508466 77698 508702 77934
rect 508466 77378 508702 77614
rect 508466 41698 508702 41934
rect 508466 41378 508702 41614
rect 508466 5698 508702 5934
rect 508466 5378 508702 5614
rect 508466 -2422 508702 -2186
rect 508466 -2742 508702 -2506
rect 511946 693178 512182 693414
rect 511946 692858 512182 693094
rect 511946 657178 512182 657414
rect 511946 656858 512182 657094
rect 511946 621178 512182 621414
rect 511946 620858 512182 621094
rect 511946 585178 512182 585414
rect 511946 584858 512182 585094
rect 511946 549178 512182 549414
rect 511946 548858 512182 549094
rect 511946 513178 512182 513414
rect 511946 512858 512182 513094
rect 511946 477178 512182 477414
rect 511946 476858 512182 477094
rect 511946 441178 512182 441414
rect 511946 440858 512182 441094
rect 511946 405178 512182 405414
rect 511946 404858 512182 405094
rect 511946 369178 512182 369414
rect 511946 368858 512182 369094
rect 511946 333178 512182 333414
rect 511946 332858 512182 333094
rect 511946 297178 512182 297414
rect 511946 296858 512182 297094
rect 511946 261178 512182 261414
rect 511946 260858 512182 261094
rect 511946 225178 512182 225414
rect 511946 224858 512182 225094
rect 511946 189178 512182 189414
rect 511946 188858 512182 189094
rect 511946 153178 512182 153414
rect 511946 152858 512182 153094
rect 511946 117178 512182 117414
rect 511946 116858 512182 117094
rect 511946 81178 512182 81414
rect 511946 80858 512182 81094
rect 511946 45178 512182 45414
rect 511946 44858 512182 45094
rect 511946 9178 512182 9414
rect 511946 8858 512182 9094
rect 511946 -4262 512182 -4026
rect 511946 -4582 512182 -4346
rect 533426 711042 533662 711278
rect 533426 710722 533662 710958
rect 529946 709202 530182 709438
rect 529946 708882 530182 709118
rect 526466 707362 526702 707598
rect 526466 707042 526702 707278
rect 515426 696658 515662 696894
rect 515426 696338 515662 696574
rect 515426 660658 515662 660894
rect 515426 660338 515662 660574
rect 515426 624658 515662 624894
rect 515426 624338 515662 624574
rect 515426 588658 515662 588894
rect 515426 588338 515662 588574
rect 515426 552658 515662 552894
rect 515426 552338 515662 552574
rect 515426 516658 515662 516894
rect 515426 516338 515662 516574
rect 515426 480658 515662 480894
rect 515426 480338 515662 480574
rect 515426 444658 515662 444894
rect 515426 444338 515662 444574
rect 515426 408658 515662 408894
rect 515426 408338 515662 408574
rect 515426 372658 515662 372894
rect 515426 372338 515662 372574
rect 515426 336658 515662 336894
rect 515426 336338 515662 336574
rect 515426 300658 515662 300894
rect 515426 300338 515662 300574
rect 515426 264658 515662 264894
rect 515426 264338 515662 264574
rect 515426 228658 515662 228894
rect 515426 228338 515662 228574
rect 515426 192658 515662 192894
rect 515426 192338 515662 192574
rect 515426 156658 515662 156894
rect 515426 156338 515662 156574
rect 515426 120658 515662 120894
rect 515426 120338 515662 120574
rect 515426 84658 515662 84894
rect 515426 84338 515662 84574
rect 515426 48658 515662 48894
rect 515426 48338 515662 48574
rect 515426 12658 515662 12894
rect 515426 12338 515662 12574
rect 497426 -7022 497662 -6786
rect 497426 -7342 497662 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526466 671698 526702 671934
rect 526466 671378 526702 671614
rect 526466 635698 526702 635934
rect 526466 635378 526702 635614
rect 526466 599698 526702 599934
rect 526466 599378 526702 599614
rect 526466 563698 526702 563934
rect 526466 563378 526702 563614
rect 526466 527698 526702 527934
rect 526466 527378 526702 527614
rect 526466 491698 526702 491934
rect 526466 491378 526702 491614
rect 526466 455698 526702 455934
rect 526466 455378 526702 455614
rect 526466 419698 526702 419934
rect 526466 419378 526702 419614
rect 526466 383698 526702 383934
rect 526466 383378 526702 383614
rect 526466 347698 526702 347934
rect 526466 347378 526702 347614
rect 526466 311698 526702 311934
rect 526466 311378 526702 311614
rect 526466 275698 526702 275934
rect 526466 275378 526702 275614
rect 526466 239698 526702 239934
rect 526466 239378 526702 239614
rect 526466 203698 526702 203934
rect 526466 203378 526702 203614
rect 526466 167698 526702 167934
rect 526466 167378 526702 167614
rect 526466 131698 526702 131934
rect 526466 131378 526702 131614
rect 526466 95698 526702 95934
rect 526466 95378 526702 95614
rect 526466 59698 526702 59934
rect 526466 59378 526702 59614
rect 526466 23698 526702 23934
rect 526466 23378 526702 23614
rect 526466 -3342 526702 -3106
rect 526466 -3662 526702 -3426
rect 529946 675178 530182 675414
rect 529946 674858 530182 675094
rect 529946 639178 530182 639414
rect 529946 638858 530182 639094
rect 529946 603178 530182 603414
rect 529946 602858 530182 603094
rect 529946 567178 530182 567414
rect 529946 566858 530182 567094
rect 529946 531178 530182 531414
rect 529946 530858 530182 531094
rect 529946 495178 530182 495414
rect 529946 494858 530182 495094
rect 529946 459178 530182 459414
rect 529946 458858 530182 459094
rect 529946 423178 530182 423414
rect 529946 422858 530182 423094
rect 529946 387178 530182 387414
rect 529946 386858 530182 387094
rect 529946 351178 530182 351414
rect 529946 350858 530182 351094
rect 529946 315178 530182 315414
rect 529946 314858 530182 315094
rect 529946 279178 530182 279414
rect 529946 278858 530182 279094
rect 529946 243178 530182 243414
rect 529946 242858 530182 243094
rect 529946 207178 530182 207414
rect 529946 206858 530182 207094
rect 529946 171178 530182 171414
rect 529946 170858 530182 171094
rect 529946 135178 530182 135414
rect 529946 134858 530182 135094
rect 529946 99178 530182 99414
rect 529946 98858 530182 99094
rect 529946 63178 530182 63414
rect 529946 62858 530182 63094
rect 529946 27178 530182 27414
rect 529946 26858 530182 27094
rect 529946 -5182 530182 -4946
rect 529946 -5502 530182 -5266
rect 551426 710122 551662 710358
rect 551426 709802 551662 710038
rect 547946 708282 548182 708518
rect 547946 707962 548182 708198
rect 544466 706442 544702 706678
rect 544466 706122 544702 706358
rect 533426 678658 533662 678894
rect 533426 678338 533662 678574
rect 533426 642658 533662 642894
rect 533426 642338 533662 642574
rect 533426 606658 533662 606894
rect 533426 606338 533662 606574
rect 533426 570658 533662 570894
rect 533426 570338 533662 570574
rect 533426 534658 533662 534894
rect 533426 534338 533662 534574
rect 533426 498658 533662 498894
rect 533426 498338 533662 498574
rect 533426 462658 533662 462894
rect 533426 462338 533662 462574
rect 533426 426658 533662 426894
rect 533426 426338 533662 426574
rect 533426 390658 533662 390894
rect 533426 390338 533662 390574
rect 533426 354658 533662 354894
rect 533426 354338 533662 354574
rect 533426 318658 533662 318894
rect 533426 318338 533662 318574
rect 533426 282658 533662 282894
rect 533426 282338 533662 282574
rect 533426 246658 533662 246894
rect 533426 246338 533662 246574
rect 533426 210658 533662 210894
rect 533426 210338 533662 210574
rect 533426 174658 533662 174894
rect 533426 174338 533662 174574
rect 533426 138658 533662 138894
rect 533426 138338 533662 138574
rect 533426 102658 533662 102894
rect 533426 102338 533662 102574
rect 533426 66658 533662 66894
rect 533426 66338 533662 66574
rect 533426 30658 533662 30894
rect 533426 30338 533662 30574
rect 515426 -6102 515662 -5866
rect 515426 -6422 515662 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544466 689698 544702 689934
rect 544466 689378 544702 689614
rect 544466 653698 544702 653934
rect 544466 653378 544702 653614
rect 544466 617698 544702 617934
rect 544466 617378 544702 617614
rect 544466 581698 544702 581934
rect 544466 581378 544702 581614
rect 544466 545698 544702 545934
rect 544466 545378 544702 545614
rect 544466 509698 544702 509934
rect 544466 509378 544702 509614
rect 544466 473698 544702 473934
rect 544466 473378 544702 473614
rect 544466 437698 544702 437934
rect 544466 437378 544702 437614
rect 544466 401698 544702 401934
rect 544466 401378 544702 401614
rect 544466 365698 544702 365934
rect 544466 365378 544702 365614
rect 544466 329698 544702 329934
rect 544466 329378 544702 329614
rect 544466 293698 544702 293934
rect 544466 293378 544702 293614
rect 544466 257698 544702 257934
rect 544466 257378 544702 257614
rect 544466 221698 544702 221934
rect 544466 221378 544702 221614
rect 544466 185698 544702 185934
rect 544466 185378 544702 185614
rect 544466 149698 544702 149934
rect 544466 149378 544702 149614
rect 544466 113698 544702 113934
rect 544466 113378 544702 113614
rect 544466 77698 544702 77934
rect 544466 77378 544702 77614
rect 544466 41698 544702 41934
rect 544466 41378 544702 41614
rect 544466 5698 544702 5934
rect 544466 5378 544702 5614
rect 544466 -2422 544702 -2186
rect 544466 -2742 544702 -2506
rect 547946 693178 548182 693414
rect 547946 692858 548182 693094
rect 547946 657178 548182 657414
rect 547946 656858 548182 657094
rect 547946 621178 548182 621414
rect 547946 620858 548182 621094
rect 547946 585178 548182 585414
rect 547946 584858 548182 585094
rect 547946 549178 548182 549414
rect 547946 548858 548182 549094
rect 547946 513178 548182 513414
rect 547946 512858 548182 513094
rect 547946 477178 548182 477414
rect 547946 476858 548182 477094
rect 547946 441178 548182 441414
rect 547946 440858 548182 441094
rect 547946 405178 548182 405414
rect 547946 404858 548182 405094
rect 547946 369178 548182 369414
rect 547946 368858 548182 369094
rect 547946 333178 548182 333414
rect 547946 332858 548182 333094
rect 547946 297178 548182 297414
rect 547946 296858 548182 297094
rect 547946 261178 548182 261414
rect 547946 260858 548182 261094
rect 547946 225178 548182 225414
rect 547946 224858 548182 225094
rect 547946 189178 548182 189414
rect 547946 188858 548182 189094
rect 547946 153178 548182 153414
rect 547946 152858 548182 153094
rect 547946 117178 548182 117414
rect 547946 116858 548182 117094
rect 547946 81178 548182 81414
rect 547946 80858 548182 81094
rect 547946 45178 548182 45414
rect 547946 44858 548182 45094
rect 547946 9178 548182 9414
rect 547946 8858 548182 9094
rect 547946 -4262 548182 -4026
rect 547946 -4582 548182 -4346
rect 569426 711042 569662 711278
rect 569426 710722 569662 710958
rect 565946 709202 566182 709438
rect 565946 708882 566182 709118
rect 562466 707362 562702 707598
rect 562466 707042 562702 707278
rect 551426 696658 551662 696894
rect 551426 696338 551662 696574
rect 551426 660658 551662 660894
rect 551426 660338 551662 660574
rect 551426 624658 551662 624894
rect 551426 624338 551662 624574
rect 551426 588658 551662 588894
rect 551426 588338 551662 588574
rect 551426 552658 551662 552894
rect 551426 552338 551662 552574
rect 551426 516658 551662 516894
rect 551426 516338 551662 516574
rect 551426 480658 551662 480894
rect 551426 480338 551662 480574
rect 551426 444658 551662 444894
rect 551426 444338 551662 444574
rect 551426 408658 551662 408894
rect 551426 408338 551662 408574
rect 551426 372658 551662 372894
rect 551426 372338 551662 372574
rect 551426 336658 551662 336894
rect 551426 336338 551662 336574
rect 551426 300658 551662 300894
rect 551426 300338 551662 300574
rect 551426 264658 551662 264894
rect 551426 264338 551662 264574
rect 551426 228658 551662 228894
rect 551426 228338 551662 228574
rect 551426 192658 551662 192894
rect 551426 192338 551662 192574
rect 551426 156658 551662 156894
rect 551426 156338 551662 156574
rect 551426 120658 551662 120894
rect 551426 120338 551662 120574
rect 551426 84658 551662 84894
rect 551426 84338 551662 84574
rect 551426 48658 551662 48894
rect 551426 48338 551662 48574
rect 551426 12658 551662 12894
rect 551426 12338 551662 12574
rect 533426 -7022 533662 -6786
rect 533426 -7342 533662 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562466 671698 562702 671934
rect 562466 671378 562702 671614
rect 562466 635698 562702 635934
rect 562466 635378 562702 635614
rect 562466 599698 562702 599934
rect 562466 599378 562702 599614
rect 562466 563698 562702 563934
rect 562466 563378 562702 563614
rect 562466 527698 562702 527934
rect 562466 527378 562702 527614
rect 562466 491698 562702 491934
rect 562466 491378 562702 491614
rect 562466 455698 562702 455934
rect 562466 455378 562702 455614
rect 562466 419698 562702 419934
rect 562466 419378 562702 419614
rect 562466 383698 562702 383934
rect 562466 383378 562702 383614
rect 562466 347698 562702 347934
rect 562466 347378 562702 347614
rect 562466 311698 562702 311934
rect 562466 311378 562702 311614
rect 562466 275698 562702 275934
rect 562466 275378 562702 275614
rect 562466 239698 562702 239934
rect 562466 239378 562702 239614
rect 562466 203698 562702 203934
rect 562466 203378 562702 203614
rect 562466 167698 562702 167934
rect 562466 167378 562702 167614
rect 562466 131698 562702 131934
rect 562466 131378 562702 131614
rect 562466 95698 562702 95934
rect 562466 95378 562702 95614
rect 562466 59698 562702 59934
rect 562466 59378 562702 59614
rect 562466 23698 562702 23934
rect 562466 23378 562702 23614
rect 562466 -3342 562702 -3106
rect 562466 -3662 562702 -3426
rect 565946 675178 566182 675414
rect 565946 674858 566182 675094
rect 565946 639178 566182 639414
rect 565946 638858 566182 639094
rect 565946 603178 566182 603414
rect 565946 602858 566182 603094
rect 565946 567178 566182 567414
rect 565946 566858 566182 567094
rect 565946 531178 566182 531414
rect 565946 530858 566182 531094
rect 565946 495178 566182 495414
rect 565946 494858 566182 495094
rect 565946 459178 566182 459414
rect 565946 458858 566182 459094
rect 565946 423178 566182 423414
rect 565946 422858 566182 423094
rect 565946 387178 566182 387414
rect 565946 386858 566182 387094
rect 565946 351178 566182 351414
rect 565946 350858 566182 351094
rect 565946 315178 566182 315414
rect 565946 314858 566182 315094
rect 565946 279178 566182 279414
rect 565946 278858 566182 279094
rect 565946 243178 566182 243414
rect 565946 242858 566182 243094
rect 565946 207178 566182 207414
rect 565946 206858 566182 207094
rect 565946 171178 566182 171414
rect 565946 170858 566182 171094
rect 565946 135178 566182 135414
rect 565946 134858 566182 135094
rect 565946 99178 566182 99414
rect 565946 98858 566182 99094
rect 565946 63178 566182 63414
rect 565946 62858 566182 63094
rect 565946 27178 566182 27414
rect 565946 26858 566182 27094
rect 565946 -5182 566182 -4946
rect 565946 -5502 566182 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580466 706442 580702 706678
rect 580466 706122 580702 706358
rect 569426 678658 569662 678894
rect 569426 678338 569662 678574
rect 569426 642658 569662 642894
rect 569426 642338 569662 642574
rect 569426 606658 569662 606894
rect 569426 606338 569662 606574
rect 569426 570658 569662 570894
rect 569426 570338 569662 570574
rect 569426 534658 569662 534894
rect 569426 534338 569662 534574
rect 569426 498658 569662 498894
rect 569426 498338 569662 498574
rect 569426 462658 569662 462894
rect 569426 462338 569662 462574
rect 569426 426658 569662 426894
rect 569426 426338 569662 426574
rect 569426 390658 569662 390894
rect 569426 390338 569662 390574
rect 569426 354658 569662 354894
rect 569426 354338 569662 354574
rect 569426 318658 569662 318894
rect 569426 318338 569662 318574
rect 569426 282658 569662 282894
rect 569426 282338 569662 282574
rect 569426 246658 569662 246894
rect 569426 246338 569662 246574
rect 569426 210658 569662 210894
rect 569426 210338 569662 210574
rect 569426 174658 569662 174894
rect 569426 174338 569662 174574
rect 569426 138658 569662 138894
rect 569426 138338 569662 138574
rect 569426 102658 569662 102894
rect 569426 102338 569662 102574
rect 569426 66658 569662 66894
rect 569426 66338 569662 66574
rect 569426 30658 569662 30894
rect 569426 30338 569662 30574
rect 551426 -6102 551662 -5866
rect 551426 -6422 551662 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580466 689698 580702 689934
rect 580466 689378 580702 689614
rect 580466 653698 580702 653934
rect 580466 653378 580702 653614
rect 580466 617698 580702 617934
rect 580466 617378 580702 617614
rect 580466 581698 580702 581934
rect 580466 581378 580702 581614
rect 580466 545698 580702 545934
rect 580466 545378 580702 545614
rect 580466 509698 580702 509934
rect 580466 509378 580702 509614
rect 580466 473698 580702 473934
rect 580466 473378 580702 473614
rect 580466 437698 580702 437934
rect 580466 437378 580702 437614
rect 580466 401698 580702 401934
rect 580466 401378 580702 401614
rect 580466 365698 580702 365934
rect 580466 365378 580702 365614
rect 580466 329698 580702 329934
rect 580466 329378 580702 329614
rect 580466 293698 580702 293934
rect 580466 293378 580702 293614
rect 580466 257698 580702 257934
rect 580466 257378 580702 257614
rect 580466 221698 580702 221934
rect 580466 221378 580702 221614
rect 580466 185698 580702 185934
rect 580466 185378 580702 185614
rect 580466 149698 580702 149934
rect 580466 149378 580702 149614
rect 580466 113698 580702 113934
rect 580466 113378 580702 113614
rect 580466 77698 580702 77934
rect 580466 77378 580702 77614
rect 580466 41698 580702 41934
rect 580466 41378 580702 41614
rect 580466 5698 580702 5934
rect 580466 5378 580702 5614
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689698 587578 689934
rect 587342 689378 587578 689614
rect 587342 653698 587578 653934
rect 587342 653378 587578 653614
rect 587342 617698 587578 617934
rect 587342 617378 587578 617614
rect 587342 581698 587578 581934
rect 587342 581378 587578 581614
rect 587342 545698 587578 545934
rect 587342 545378 587578 545614
rect 587342 509698 587578 509934
rect 587342 509378 587578 509614
rect 587342 473698 587578 473934
rect 587342 473378 587578 473614
rect 587342 437698 587578 437934
rect 587342 437378 587578 437614
rect 587342 401698 587578 401934
rect 587342 401378 587578 401614
rect 587342 365698 587578 365934
rect 587342 365378 587578 365614
rect 587342 329698 587578 329934
rect 587342 329378 587578 329614
rect 587342 293698 587578 293934
rect 587342 293378 587578 293614
rect 587342 257698 587578 257934
rect 587342 257378 587578 257614
rect 587342 221698 587578 221934
rect 587342 221378 587578 221614
rect 587342 185698 587578 185934
rect 587342 185378 587578 185614
rect 587342 149698 587578 149934
rect 587342 149378 587578 149614
rect 587342 113698 587578 113934
rect 587342 113378 587578 113614
rect 587342 77698 587578 77934
rect 587342 77378 587578 77614
rect 587342 41698 587578 41934
rect 587342 41378 587578 41614
rect 587342 5698 587578 5934
rect 587342 5378 587578 5614
rect 580466 -2422 580702 -2186
rect 580466 -2742 580702 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671698 588498 671934
rect 588262 671378 588498 671614
rect 588262 635698 588498 635934
rect 588262 635378 588498 635614
rect 588262 599698 588498 599934
rect 588262 599378 588498 599614
rect 588262 563698 588498 563934
rect 588262 563378 588498 563614
rect 588262 527698 588498 527934
rect 588262 527378 588498 527614
rect 588262 491698 588498 491934
rect 588262 491378 588498 491614
rect 588262 455698 588498 455934
rect 588262 455378 588498 455614
rect 588262 419698 588498 419934
rect 588262 419378 588498 419614
rect 588262 383698 588498 383934
rect 588262 383378 588498 383614
rect 588262 347698 588498 347934
rect 588262 347378 588498 347614
rect 588262 311698 588498 311934
rect 588262 311378 588498 311614
rect 588262 275698 588498 275934
rect 588262 275378 588498 275614
rect 588262 239698 588498 239934
rect 588262 239378 588498 239614
rect 588262 203698 588498 203934
rect 588262 203378 588498 203614
rect 588262 167698 588498 167934
rect 588262 167378 588498 167614
rect 588262 131698 588498 131934
rect 588262 131378 588498 131614
rect 588262 95698 588498 95934
rect 588262 95378 588498 95614
rect 588262 59698 588498 59934
rect 588262 59378 588498 59614
rect 588262 23698 588498 23934
rect 588262 23378 588498 23614
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693178 589418 693414
rect 589182 692858 589418 693094
rect 589182 657178 589418 657414
rect 589182 656858 589418 657094
rect 589182 621178 589418 621414
rect 589182 620858 589418 621094
rect 589182 585178 589418 585414
rect 589182 584858 589418 585094
rect 589182 549178 589418 549414
rect 589182 548858 589418 549094
rect 589182 513178 589418 513414
rect 589182 512858 589418 513094
rect 589182 477178 589418 477414
rect 589182 476858 589418 477094
rect 589182 441178 589418 441414
rect 589182 440858 589418 441094
rect 589182 405178 589418 405414
rect 589182 404858 589418 405094
rect 589182 369178 589418 369414
rect 589182 368858 589418 369094
rect 589182 333178 589418 333414
rect 589182 332858 589418 333094
rect 589182 297178 589418 297414
rect 589182 296858 589418 297094
rect 589182 261178 589418 261414
rect 589182 260858 589418 261094
rect 589182 225178 589418 225414
rect 589182 224858 589418 225094
rect 589182 189178 589418 189414
rect 589182 188858 589418 189094
rect 589182 153178 589418 153414
rect 589182 152858 589418 153094
rect 589182 117178 589418 117414
rect 589182 116858 589418 117094
rect 589182 81178 589418 81414
rect 589182 80858 589418 81094
rect 589182 45178 589418 45414
rect 589182 44858 589418 45094
rect 589182 9178 589418 9414
rect 589182 8858 589418 9094
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675178 590338 675414
rect 590102 674858 590338 675094
rect 590102 639178 590338 639414
rect 590102 638858 590338 639094
rect 590102 603178 590338 603414
rect 590102 602858 590338 603094
rect 590102 567178 590338 567414
rect 590102 566858 590338 567094
rect 590102 531178 590338 531414
rect 590102 530858 590338 531094
rect 590102 495178 590338 495414
rect 590102 494858 590338 495094
rect 590102 459178 590338 459414
rect 590102 458858 590338 459094
rect 590102 423178 590338 423414
rect 590102 422858 590338 423094
rect 590102 387178 590338 387414
rect 590102 386858 590338 387094
rect 590102 351178 590338 351414
rect 590102 350858 590338 351094
rect 590102 315178 590338 315414
rect 590102 314858 590338 315094
rect 590102 279178 590338 279414
rect 590102 278858 590338 279094
rect 590102 243178 590338 243414
rect 590102 242858 590338 243094
rect 590102 207178 590338 207414
rect 590102 206858 590338 207094
rect 590102 171178 590338 171414
rect 590102 170858 590338 171094
rect 590102 135178 590338 135414
rect 590102 134858 590338 135094
rect 590102 99178 590338 99414
rect 590102 98858 590338 99094
rect 590102 63178 590338 63414
rect 590102 62858 590338 63094
rect 590102 27178 590338 27414
rect 590102 26858 590338 27094
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 696658 591258 696894
rect 591022 696338 591258 696574
rect 591022 660658 591258 660894
rect 591022 660338 591258 660574
rect 591022 624658 591258 624894
rect 591022 624338 591258 624574
rect 591022 588658 591258 588894
rect 591022 588338 591258 588574
rect 591022 552658 591258 552894
rect 591022 552338 591258 552574
rect 591022 516658 591258 516894
rect 591022 516338 591258 516574
rect 591022 480658 591258 480894
rect 591022 480338 591258 480574
rect 591022 444658 591258 444894
rect 591022 444338 591258 444574
rect 591022 408658 591258 408894
rect 591022 408338 591258 408574
rect 591022 372658 591258 372894
rect 591022 372338 591258 372574
rect 591022 336658 591258 336894
rect 591022 336338 591258 336574
rect 591022 300658 591258 300894
rect 591022 300338 591258 300574
rect 591022 264658 591258 264894
rect 591022 264338 591258 264574
rect 591022 228658 591258 228894
rect 591022 228338 591258 228574
rect 591022 192658 591258 192894
rect 591022 192338 591258 192574
rect 591022 156658 591258 156894
rect 591022 156338 591258 156574
rect 591022 120658 591258 120894
rect 591022 120338 591258 120574
rect 591022 84658 591258 84894
rect 591022 84338 591258 84574
rect 591022 48658 591258 48894
rect 591022 48338 591258 48574
rect 591022 12658 591258 12894
rect 591022 12338 591258 12574
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 678658 592178 678894
rect 591942 678338 592178 678574
rect 591942 642658 592178 642894
rect 591942 642338 592178 642574
rect 591942 606658 592178 606894
rect 591942 606338 592178 606574
rect 591942 570658 592178 570894
rect 591942 570338 592178 570574
rect 591942 534658 592178 534894
rect 591942 534338 592178 534574
rect 591942 498658 592178 498894
rect 591942 498338 592178 498574
rect 591942 462658 592178 462894
rect 591942 462338 592178 462574
rect 591942 426658 592178 426894
rect 591942 426338 592178 426574
rect 591942 390658 592178 390894
rect 591942 390338 592178 390574
rect 591942 354658 592178 354894
rect 591942 354338 592178 354574
rect 591942 318658 592178 318894
rect 591942 318338 592178 318574
rect 591942 282658 592178 282894
rect 591942 282338 592178 282574
rect 591942 246658 592178 246894
rect 591942 246338 592178 246574
rect 591942 210658 592178 210894
rect 591942 210338 592178 210574
rect 591942 174658 592178 174894
rect 591942 174338 592178 174574
rect 591942 138658 592178 138894
rect 591942 138338 592178 138574
rect 591942 102658 592178 102894
rect 591942 102338 592178 102574
rect 591942 66658 592178 66894
rect 591942 66338 592178 66574
rect 591942 30658 592178 30894
rect 591942 30338 592178 30574
rect 569426 -7022 569662 -6786
rect 569426 -7342 569662 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8426 711290 -7846 711302
rect 29254 711290 29834 711302
rect 65254 711290 65834 711302
rect 101254 711290 101834 711302
rect 137254 711290 137834 711302
rect 173254 711290 173834 711302
rect 209254 711290 209834 711302
rect 245254 711290 245834 711302
rect 281254 711290 281834 711302
rect 317254 711290 317834 711302
rect 353254 711290 353834 711302
rect 389254 711290 389834 711302
rect 425254 711290 425834 711302
rect 461254 711290 461834 711302
rect 497254 711290 497834 711302
rect 533254 711290 533834 711302
rect 569254 711290 569834 711302
rect 591770 711290 592350 711302
rect -8426 711278 592350 711290
rect -8426 711042 -8254 711278
rect -8018 711042 29426 711278
rect 29662 711042 65426 711278
rect 65662 711042 101426 711278
rect 101662 711042 137426 711278
rect 137662 711042 173426 711278
rect 173662 711042 209426 711278
rect 209662 711042 245426 711278
rect 245662 711042 281426 711278
rect 281662 711042 317426 711278
rect 317662 711042 353426 711278
rect 353662 711042 389426 711278
rect 389662 711042 425426 711278
rect 425662 711042 461426 711278
rect 461662 711042 497426 711278
rect 497662 711042 533426 711278
rect 533662 711042 569426 711278
rect 569662 711042 591942 711278
rect 592178 711042 592350 711278
rect -8426 710958 592350 711042
rect -8426 710722 -8254 710958
rect -8018 710722 29426 710958
rect 29662 710722 65426 710958
rect 65662 710722 101426 710958
rect 101662 710722 137426 710958
rect 137662 710722 173426 710958
rect 173662 710722 209426 710958
rect 209662 710722 245426 710958
rect 245662 710722 281426 710958
rect 281662 710722 317426 710958
rect 317662 710722 353426 710958
rect 353662 710722 389426 710958
rect 389662 710722 425426 710958
rect 425662 710722 461426 710958
rect 461662 710722 497426 710958
rect 497662 710722 533426 710958
rect 533662 710722 569426 710958
rect 569662 710722 591942 710958
rect 592178 710722 592350 710958
rect -8426 710710 592350 710722
rect -8426 710698 -7846 710710
rect 29254 710698 29834 710710
rect 65254 710698 65834 710710
rect 101254 710698 101834 710710
rect 137254 710698 137834 710710
rect 173254 710698 173834 710710
rect 209254 710698 209834 710710
rect 245254 710698 245834 710710
rect 281254 710698 281834 710710
rect 317254 710698 317834 710710
rect 353254 710698 353834 710710
rect 389254 710698 389834 710710
rect 425254 710698 425834 710710
rect 461254 710698 461834 710710
rect 497254 710698 497834 710710
rect 533254 710698 533834 710710
rect 569254 710698 569834 710710
rect 591770 710698 592350 710710
rect -7506 710370 -6926 710382
rect 11254 710370 11834 710382
rect 47254 710370 47834 710382
rect 83254 710370 83834 710382
rect 119254 710370 119834 710382
rect 155254 710370 155834 710382
rect 191254 710370 191834 710382
rect 227254 710370 227834 710382
rect 263254 710370 263834 710382
rect 299254 710370 299834 710382
rect 335254 710370 335834 710382
rect 371254 710370 371834 710382
rect 407254 710370 407834 710382
rect 443254 710370 443834 710382
rect 479254 710370 479834 710382
rect 515254 710370 515834 710382
rect 551254 710370 551834 710382
rect 590850 710370 591430 710382
rect -7506 710358 591430 710370
rect -7506 710122 -7334 710358
rect -7098 710122 11426 710358
rect 11662 710122 47426 710358
rect 47662 710122 83426 710358
rect 83662 710122 119426 710358
rect 119662 710122 155426 710358
rect 155662 710122 191426 710358
rect 191662 710122 227426 710358
rect 227662 710122 263426 710358
rect 263662 710122 299426 710358
rect 299662 710122 335426 710358
rect 335662 710122 371426 710358
rect 371662 710122 407426 710358
rect 407662 710122 443426 710358
rect 443662 710122 479426 710358
rect 479662 710122 515426 710358
rect 515662 710122 551426 710358
rect 551662 710122 591022 710358
rect 591258 710122 591430 710358
rect -7506 710038 591430 710122
rect -7506 709802 -7334 710038
rect -7098 709802 11426 710038
rect 11662 709802 47426 710038
rect 47662 709802 83426 710038
rect 83662 709802 119426 710038
rect 119662 709802 155426 710038
rect 155662 709802 191426 710038
rect 191662 709802 227426 710038
rect 227662 709802 263426 710038
rect 263662 709802 299426 710038
rect 299662 709802 335426 710038
rect 335662 709802 371426 710038
rect 371662 709802 407426 710038
rect 407662 709802 443426 710038
rect 443662 709802 479426 710038
rect 479662 709802 515426 710038
rect 515662 709802 551426 710038
rect 551662 709802 591022 710038
rect 591258 709802 591430 710038
rect -7506 709790 591430 709802
rect -7506 709778 -6926 709790
rect 11254 709778 11834 709790
rect 47254 709778 47834 709790
rect 83254 709778 83834 709790
rect 119254 709778 119834 709790
rect 155254 709778 155834 709790
rect 191254 709778 191834 709790
rect 227254 709778 227834 709790
rect 263254 709778 263834 709790
rect 299254 709778 299834 709790
rect 335254 709778 335834 709790
rect 371254 709778 371834 709790
rect 407254 709778 407834 709790
rect 443254 709778 443834 709790
rect 479254 709778 479834 709790
rect 515254 709778 515834 709790
rect 551254 709778 551834 709790
rect 590850 709778 591430 709790
rect -6586 709450 -6006 709462
rect 25774 709450 26354 709462
rect 61774 709450 62354 709462
rect 97774 709450 98354 709462
rect 133774 709450 134354 709462
rect 169774 709450 170354 709462
rect 205774 709450 206354 709462
rect 241774 709450 242354 709462
rect 277774 709450 278354 709462
rect 313774 709450 314354 709462
rect 349774 709450 350354 709462
rect 385774 709450 386354 709462
rect 421774 709450 422354 709462
rect 457774 709450 458354 709462
rect 493774 709450 494354 709462
rect 529774 709450 530354 709462
rect 565774 709450 566354 709462
rect 589930 709450 590510 709462
rect -6586 709438 590510 709450
rect -6586 709202 -6414 709438
rect -6178 709202 25946 709438
rect 26182 709202 61946 709438
rect 62182 709202 97946 709438
rect 98182 709202 133946 709438
rect 134182 709202 169946 709438
rect 170182 709202 205946 709438
rect 206182 709202 241946 709438
rect 242182 709202 277946 709438
rect 278182 709202 313946 709438
rect 314182 709202 349946 709438
rect 350182 709202 385946 709438
rect 386182 709202 421946 709438
rect 422182 709202 457946 709438
rect 458182 709202 493946 709438
rect 494182 709202 529946 709438
rect 530182 709202 565946 709438
rect 566182 709202 590102 709438
rect 590338 709202 590510 709438
rect -6586 709118 590510 709202
rect -6586 708882 -6414 709118
rect -6178 708882 25946 709118
rect 26182 708882 61946 709118
rect 62182 708882 97946 709118
rect 98182 708882 133946 709118
rect 134182 708882 169946 709118
rect 170182 708882 205946 709118
rect 206182 708882 241946 709118
rect 242182 708882 277946 709118
rect 278182 708882 313946 709118
rect 314182 708882 349946 709118
rect 350182 708882 385946 709118
rect 386182 708882 421946 709118
rect 422182 708882 457946 709118
rect 458182 708882 493946 709118
rect 494182 708882 529946 709118
rect 530182 708882 565946 709118
rect 566182 708882 590102 709118
rect 590338 708882 590510 709118
rect -6586 708870 590510 708882
rect -6586 708858 -6006 708870
rect 25774 708858 26354 708870
rect 61774 708858 62354 708870
rect 97774 708858 98354 708870
rect 133774 708858 134354 708870
rect 169774 708858 170354 708870
rect 205774 708858 206354 708870
rect 241774 708858 242354 708870
rect 277774 708858 278354 708870
rect 313774 708858 314354 708870
rect 349774 708858 350354 708870
rect 385774 708858 386354 708870
rect 421774 708858 422354 708870
rect 457774 708858 458354 708870
rect 493774 708858 494354 708870
rect 529774 708858 530354 708870
rect 565774 708858 566354 708870
rect 589930 708858 590510 708870
rect -5666 708530 -5086 708542
rect 7774 708530 8354 708542
rect 43774 708530 44354 708542
rect 79774 708530 80354 708542
rect 115774 708530 116354 708542
rect 151774 708530 152354 708542
rect 187774 708530 188354 708542
rect 223774 708530 224354 708542
rect 259774 708530 260354 708542
rect 295774 708530 296354 708542
rect 331774 708530 332354 708542
rect 367774 708530 368354 708542
rect 403774 708530 404354 708542
rect 439774 708530 440354 708542
rect 475774 708530 476354 708542
rect 511774 708530 512354 708542
rect 547774 708530 548354 708542
rect 589010 708530 589590 708542
rect -5666 708518 589590 708530
rect -5666 708282 -5494 708518
rect -5258 708282 7946 708518
rect 8182 708282 43946 708518
rect 44182 708282 79946 708518
rect 80182 708282 115946 708518
rect 116182 708282 151946 708518
rect 152182 708282 187946 708518
rect 188182 708282 223946 708518
rect 224182 708282 259946 708518
rect 260182 708282 295946 708518
rect 296182 708282 331946 708518
rect 332182 708282 367946 708518
rect 368182 708282 403946 708518
rect 404182 708282 439946 708518
rect 440182 708282 475946 708518
rect 476182 708282 511946 708518
rect 512182 708282 547946 708518
rect 548182 708282 589182 708518
rect 589418 708282 589590 708518
rect -5666 708198 589590 708282
rect -5666 707962 -5494 708198
rect -5258 707962 7946 708198
rect 8182 707962 43946 708198
rect 44182 707962 79946 708198
rect 80182 707962 115946 708198
rect 116182 707962 151946 708198
rect 152182 707962 187946 708198
rect 188182 707962 223946 708198
rect 224182 707962 259946 708198
rect 260182 707962 295946 708198
rect 296182 707962 331946 708198
rect 332182 707962 367946 708198
rect 368182 707962 403946 708198
rect 404182 707962 439946 708198
rect 440182 707962 475946 708198
rect 476182 707962 511946 708198
rect 512182 707962 547946 708198
rect 548182 707962 589182 708198
rect 589418 707962 589590 708198
rect -5666 707950 589590 707962
rect -5666 707938 -5086 707950
rect 7774 707938 8354 707950
rect 43774 707938 44354 707950
rect 79774 707938 80354 707950
rect 115774 707938 116354 707950
rect 151774 707938 152354 707950
rect 187774 707938 188354 707950
rect 223774 707938 224354 707950
rect 259774 707938 260354 707950
rect 295774 707938 296354 707950
rect 331774 707938 332354 707950
rect 367774 707938 368354 707950
rect 403774 707938 404354 707950
rect 439774 707938 440354 707950
rect 475774 707938 476354 707950
rect 511774 707938 512354 707950
rect 547774 707938 548354 707950
rect 589010 707938 589590 707950
rect -4746 707610 -4166 707622
rect 22294 707610 22874 707622
rect 58294 707610 58874 707622
rect 94294 707610 94874 707622
rect 130294 707610 130874 707622
rect 166294 707610 166874 707622
rect 202294 707610 202874 707622
rect 238294 707610 238874 707622
rect 274294 707610 274874 707622
rect 310294 707610 310874 707622
rect 346294 707610 346874 707622
rect 382294 707610 382874 707622
rect 418294 707610 418874 707622
rect 454294 707610 454874 707622
rect 490294 707610 490874 707622
rect 526294 707610 526874 707622
rect 562294 707610 562874 707622
rect 588090 707610 588670 707622
rect -4746 707598 588670 707610
rect -4746 707362 -4574 707598
rect -4338 707362 22466 707598
rect 22702 707362 58466 707598
rect 58702 707362 94466 707598
rect 94702 707362 130466 707598
rect 130702 707362 166466 707598
rect 166702 707362 202466 707598
rect 202702 707362 238466 707598
rect 238702 707362 274466 707598
rect 274702 707362 310466 707598
rect 310702 707362 346466 707598
rect 346702 707362 382466 707598
rect 382702 707362 418466 707598
rect 418702 707362 454466 707598
rect 454702 707362 490466 707598
rect 490702 707362 526466 707598
rect 526702 707362 562466 707598
rect 562702 707362 588262 707598
rect 588498 707362 588670 707598
rect -4746 707278 588670 707362
rect -4746 707042 -4574 707278
rect -4338 707042 22466 707278
rect 22702 707042 58466 707278
rect 58702 707042 94466 707278
rect 94702 707042 130466 707278
rect 130702 707042 166466 707278
rect 166702 707042 202466 707278
rect 202702 707042 238466 707278
rect 238702 707042 274466 707278
rect 274702 707042 310466 707278
rect 310702 707042 346466 707278
rect 346702 707042 382466 707278
rect 382702 707042 418466 707278
rect 418702 707042 454466 707278
rect 454702 707042 490466 707278
rect 490702 707042 526466 707278
rect 526702 707042 562466 707278
rect 562702 707042 588262 707278
rect 588498 707042 588670 707278
rect -4746 707030 588670 707042
rect -4746 707018 -4166 707030
rect 22294 707018 22874 707030
rect 58294 707018 58874 707030
rect 94294 707018 94874 707030
rect 130294 707018 130874 707030
rect 166294 707018 166874 707030
rect 202294 707018 202874 707030
rect 238294 707018 238874 707030
rect 274294 707018 274874 707030
rect 310294 707018 310874 707030
rect 346294 707018 346874 707030
rect 382294 707018 382874 707030
rect 418294 707018 418874 707030
rect 454294 707018 454874 707030
rect 490294 707018 490874 707030
rect 526294 707018 526874 707030
rect 562294 707018 562874 707030
rect 588090 707018 588670 707030
rect -3826 706690 -3246 706702
rect 4294 706690 4874 706702
rect 40294 706690 40874 706702
rect 76294 706690 76874 706702
rect 112294 706690 112874 706702
rect 148294 706690 148874 706702
rect 184294 706690 184874 706702
rect 220294 706690 220874 706702
rect 256294 706690 256874 706702
rect 292294 706690 292874 706702
rect 328294 706690 328874 706702
rect 364294 706690 364874 706702
rect 400294 706690 400874 706702
rect 436294 706690 436874 706702
rect 472294 706690 472874 706702
rect 508294 706690 508874 706702
rect 544294 706690 544874 706702
rect 580294 706690 580874 706702
rect 587170 706690 587750 706702
rect -3826 706678 587750 706690
rect -3826 706442 -3654 706678
rect -3418 706442 4466 706678
rect 4702 706442 40466 706678
rect 40702 706442 76466 706678
rect 76702 706442 112466 706678
rect 112702 706442 148466 706678
rect 148702 706442 184466 706678
rect 184702 706442 220466 706678
rect 220702 706442 256466 706678
rect 256702 706442 292466 706678
rect 292702 706442 328466 706678
rect 328702 706442 364466 706678
rect 364702 706442 400466 706678
rect 400702 706442 436466 706678
rect 436702 706442 472466 706678
rect 472702 706442 508466 706678
rect 508702 706442 544466 706678
rect 544702 706442 580466 706678
rect 580702 706442 587342 706678
rect 587578 706442 587750 706678
rect -3826 706358 587750 706442
rect -3826 706122 -3654 706358
rect -3418 706122 4466 706358
rect 4702 706122 40466 706358
rect 40702 706122 76466 706358
rect 76702 706122 112466 706358
rect 112702 706122 148466 706358
rect 148702 706122 184466 706358
rect 184702 706122 220466 706358
rect 220702 706122 256466 706358
rect 256702 706122 292466 706358
rect 292702 706122 328466 706358
rect 328702 706122 364466 706358
rect 364702 706122 400466 706358
rect 400702 706122 436466 706358
rect 436702 706122 472466 706358
rect 472702 706122 508466 706358
rect 508702 706122 544466 706358
rect 544702 706122 580466 706358
rect 580702 706122 587342 706358
rect 587578 706122 587750 706358
rect -3826 706110 587750 706122
rect -3826 706098 -3246 706110
rect 4294 706098 4874 706110
rect 40294 706098 40874 706110
rect 76294 706098 76874 706110
rect 112294 706098 112874 706110
rect 148294 706098 148874 706110
rect 184294 706098 184874 706110
rect 220294 706098 220874 706110
rect 256294 706098 256874 706110
rect 292294 706098 292874 706110
rect 328294 706098 328874 706110
rect 364294 706098 364874 706110
rect 400294 706098 400874 706110
rect 436294 706098 436874 706110
rect 472294 706098 472874 706110
rect 508294 706098 508874 706110
rect 544294 706098 544874 706110
rect 580294 706098 580874 706110
rect 587170 706098 587750 706110
rect -2906 705770 -2326 705782
rect 18814 705770 19394 705782
rect 54814 705770 55394 705782
rect 90814 705770 91394 705782
rect 126814 705770 127394 705782
rect 162814 705770 163394 705782
rect 198814 705770 199394 705782
rect 234814 705770 235394 705782
rect 270814 705770 271394 705782
rect 306814 705770 307394 705782
rect 342814 705770 343394 705782
rect 378814 705770 379394 705782
rect 414814 705770 415394 705782
rect 450814 705770 451394 705782
rect 486814 705770 487394 705782
rect 522814 705770 523394 705782
rect 558814 705770 559394 705782
rect 586250 705770 586830 705782
rect -2906 705758 586830 705770
rect -2906 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586830 705758
rect -2906 705438 586830 705522
rect -2906 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586830 705438
rect -2906 705190 586830 705202
rect -2906 705178 -2326 705190
rect 18814 705178 19394 705190
rect 54814 705178 55394 705190
rect 90814 705178 91394 705190
rect 126814 705178 127394 705190
rect 162814 705178 163394 705190
rect 198814 705178 199394 705190
rect 234814 705178 235394 705190
rect 270814 705178 271394 705190
rect 306814 705178 307394 705190
rect 342814 705178 343394 705190
rect 378814 705178 379394 705190
rect 414814 705178 415394 705190
rect 450814 705178 451394 705190
rect 486814 705178 487394 705190
rect 522814 705178 523394 705190
rect 558814 705178 559394 705190
rect 586250 705178 586830 705190
rect -1986 704850 -1406 704862
rect 814 704850 1394 704862
rect 36814 704850 37394 704862
rect 72814 704850 73394 704862
rect 108814 704850 109394 704862
rect 144814 704850 145394 704862
rect 180814 704850 181394 704862
rect 216814 704850 217394 704862
rect 252814 704850 253394 704862
rect 288814 704850 289394 704862
rect 324814 704850 325394 704862
rect 360814 704850 361394 704862
rect 396814 704850 397394 704862
rect 432814 704850 433394 704862
rect 468814 704850 469394 704862
rect 504814 704850 505394 704862
rect 540814 704850 541394 704862
rect 576814 704850 577394 704862
rect 585330 704850 585910 704862
rect -1986 704838 585910 704850
rect -1986 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585910 704838
rect -1986 704518 585910 704602
rect -1986 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585910 704518
rect -1986 704270 585910 704282
rect -1986 704258 -1406 704270
rect 814 704258 1394 704270
rect 36814 704258 37394 704270
rect 72814 704258 73394 704270
rect 108814 704258 109394 704270
rect 144814 704258 145394 704270
rect 180814 704258 181394 704270
rect 216814 704258 217394 704270
rect 252814 704258 253394 704270
rect 288814 704258 289394 704270
rect 324814 704258 325394 704270
rect 360814 704258 361394 704270
rect 396814 704258 397394 704270
rect 432814 704258 433394 704270
rect 468814 704258 469394 704270
rect 504814 704258 505394 704270
rect 540814 704258 541394 704270
rect 576814 704258 577394 704270
rect 585330 704258 585910 704270
rect -7506 696906 -6926 696918
rect 11254 696906 11834 696918
rect 47254 696906 47834 696918
rect 83254 696906 83834 696918
rect 119254 696906 119834 696918
rect 155254 696906 155834 696918
rect 191254 696906 191834 696918
rect 227254 696906 227834 696918
rect 263254 696906 263834 696918
rect 299254 696906 299834 696918
rect 335254 696906 335834 696918
rect 371254 696906 371834 696918
rect 407254 696906 407834 696918
rect 443254 696906 443834 696918
rect 479254 696906 479834 696918
rect 515254 696906 515834 696918
rect 551254 696906 551834 696918
rect 590850 696906 591430 696918
rect -8426 696894 592350 696906
rect -8426 696658 -7334 696894
rect -7098 696658 11426 696894
rect 11662 696658 47426 696894
rect 47662 696658 83426 696894
rect 83662 696658 119426 696894
rect 119662 696658 155426 696894
rect 155662 696658 191426 696894
rect 191662 696658 227426 696894
rect 227662 696658 263426 696894
rect 263662 696658 299426 696894
rect 299662 696658 335426 696894
rect 335662 696658 371426 696894
rect 371662 696658 407426 696894
rect 407662 696658 443426 696894
rect 443662 696658 479426 696894
rect 479662 696658 515426 696894
rect 515662 696658 551426 696894
rect 551662 696658 591022 696894
rect 591258 696658 592350 696894
rect -8426 696574 592350 696658
rect -8426 696338 -7334 696574
rect -7098 696338 11426 696574
rect 11662 696338 47426 696574
rect 47662 696338 83426 696574
rect 83662 696338 119426 696574
rect 119662 696338 155426 696574
rect 155662 696338 191426 696574
rect 191662 696338 227426 696574
rect 227662 696338 263426 696574
rect 263662 696338 299426 696574
rect 299662 696338 335426 696574
rect 335662 696338 371426 696574
rect 371662 696338 407426 696574
rect 407662 696338 443426 696574
rect 443662 696338 479426 696574
rect 479662 696338 515426 696574
rect 515662 696338 551426 696574
rect 551662 696338 591022 696574
rect 591258 696338 592350 696574
rect -8426 696326 592350 696338
rect -7506 696314 -6926 696326
rect 11254 696314 11834 696326
rect 47254 696314 47834 696326
rect 83254 696314 83834 696326
rect 119254 696314 119834 696326
rect 155254 696314 155834 696326
rect 191254 696314 191834 696326
rect 227254 696314 227834 696326
rect 263254 696314 263834 696326
rect 299254 696314 299834 696326
rect 335254 696314 335834 696326
rect 371254 696314 371834 696326
rect 407254 696314 407834 696326
rect 443254 696314 443834 696326
rect 479254 696314 479834 696326
rect 515254 696314 515834 696326
rect 551254 696314 551834 696326
rect 590850 696314 591430 696326
rect -5666 693426 -5086 693438
rect 7774 693426 8354 693438
rect 43774 693426 44354 693438
rect 79774 693426 80354 693438
rect 115774 693426 116354 693438
rect 151774 693426 152354 693438
rect 187774 693426 188354 693438
rect 223774 693426 224354 693438
rect 259774 693426 260354 693438
rect 295774 693426 296354 693438
rect 331774 693426 332354 693438
rect 367774 693426 368354 693438
rect 403774 693426 404354 693438
rect 439774 693426 440354 693438
rect 475774 693426 476354 693438
rect 511774 693426 512354 693438
rect 547774 693426 548354 693438
rect 589010 693426 589590 693438
rect -6586 693414 590510 693426
rect -6586 693178 -5494 693414
rect -5258 693178 7946 693414
rect 8182 693178 43946 693414
rect 44182 693178 79946 693414
rect 80182 693178 115946 693414
rect 116182 693178 151946 693414
rect 152182 693178 187946 693414
rect 188182 693178 223946 693414
rect 224182 693178 259946 693414
rect 260182 693178 295946 693414
rect 296182 693178 331946 693414
rect 332182 693178 367946 693414
rect 368182 693178 403946 693414
rect 404182 693178 439946 693414
rect 440182 693178 475946 693414
rect 476182 693178 511946 693414
rect 512182 693178 547946 693414
rect 548182 693178 589182 693414
rect 589418 693178 590510 693414
rect -6586 693094 590510 693178
rect -6586 692858 -5494 693094
rect -5258 692858 7946 693094
rect 8182 692858 43946 693094
rect 44182 692858 79946 693094
rect 80182 692858 115946 693094
rect 116182 692858 151946 693094
rect 152182 692858 187946 693094
rect 188182 692858 223946 693094
rect 224182 692858 259946 693094
rect 260182 692858 295946 693094
rect 296182 692858 331946 693094
rect 332182 692858 367946 693094
rect 368182 692858 403946 693094
rect 404182 692858 439946 693094
rect 440182 692858 475946 693094
rect 476182 692858 511946 693094
rect 512182 692858 547946 693094
rect 548182 692858 589182 693094
rect 589418 692858 590510 693094
rect -6586 692846 590510 692858
rect -5666 692834 -5086 692846
rect 7774 692834 8354 692846
rect 43774 692834 44354 692846
rect 79774 692834 80354 692846
rect 115774 692834 116354 692846
rect 151774 692834 152354 692846
rect 187774 692834 188354 692846
rect 223774 692834 224354 692846
rect 259774 692834 260354 692846
rect 295774 692834 296354 692846
rect 331774 692834 332354 692846
rect 367774 692834 368354 692846
rect 403774 692834 404354 692846
rect 439774 692834 440354 692846
rect 475774 692834 476354 692846
rect 511774 692834 512354 692846
rect 547774 692834 548354 692846
rect 589010 692834 589590 692846
rect -3826 689946 -3246 689958
rect 4294 689946 4874 689958
rect 40294 689946 40874 689958
rect 76294 689946 76874 689958
rect 112294 689946 112874 689958
rect 148294 689946 148874 689958
rect 184294 689946 184874 689958
rect 220294 689946 220874 689958
rect 256294 689946 256874 689958
rect 292294 689946 292874 689958
rect 328294 689946 328874 689958
rect 364294 689946 364874 689958
rect 400294 689946 400874 689958
rect 436294 689946 436874 689958
rect 472294 689946 472874 689958
rect 508294 689946 508874 689958
rect 544294 689946 544874 689958
rect 580294 689946 580874 689958
rect 587170 689946 587750 689958
rect -4746 689934 588670 689946
rect -4746 689698 -3654 689934
rect -3418 689698 4466 689934
rect 4702 689698 40466 689934
rect 40702 689698 76466 689934
rect 76702 689698 112466 689934
rect 112702 689698 148466 689934
rect 148702 689698 184466 689934
rect 184702 689698 220466 689934
rect 220702 689698 256466 689934
rect 256702 689698 292466 689934
rect 292702 689698 328466 689934
rect 328702 689698 364466 689934
rect 364702 689698 400466 689934
rect 400702 689698 436466 689934
rect 436702 689698 472466 689934
rect 472702 689698 508466 689934
rect 508702 689698 544466 689934
rect 544702 689698 580466 689934
rect 580702 689698 587342 689934
rect 587578 689698 588670 689934
rect -4746 689614 588670 689698
rect -4746 689378 -3654 689614
rect -3418 689378 4466 689614
rect 4702 689378 40466 689614
rect 40702 689378 76466 689614
rect 76702 689378 112466 689614
rect 112702 689378 148466 689614
rect 148702 689378 184466 689614
rect 184702 689378 220466 689614
rect 220702 689378 256466 689614
rect 256702 689378 292466 689614
rect 292702 689378 328466 689614
rect 328702 689378 364466 689614
rect 364702 689378 400466 689614
rect 400702 689378 436466 689614
rect 436702 689378 472466 689614
rect 472702 689378 508466 689614
rect 508702 689378 544466 689614
rect 544702 689378 580466 689614
rect 580702 689378 587342 689614
rect 587578 689378 588670 689614
rect -4746 689366 588670 689378
rect -3826 689354 -3246 689366
rect 4294 689354 4874 689366
rect 40294 689354 40874 689366
rect 76294 689354 76874 689366
rect 112294 689354 112874 689366
rect 148294 689354 148874 689366
rect 184294 689354 184874 689366
rect 220294 689354 220874 689366
rect 256294 689354 256874 689366
rect 292294 689354 292874 689366
rect 328294 689354 328874 689366
rect 364294 689354 364874 689366
rect 400294 689354 400874 689366
rect 436294 689354 436874 689366
rect 472294 689354 472874 689366
rect 508294 689354 508874 689366
rect 544294 689354 544874 689366
rect 580294 689354 580874 689366
rect 587170 689354 587750 689366
rect -1986 686466 -1406 686478
rect 814 686466 1394 686478
rect 36814 686466 37394 686478
rect 72814 686466 73394 686478
rect 108814 686466 109394 686478
rect 144814 686466 145394 686478
rect 180814 686466 181394 686478
rect 216814 686466 217394 686478
rect 252814 686466 253394 686478
rect 288814 686466 289394 686478
rect 324814 686466 325394 686478
rect 360814 686466 361394 686478
rect 396814 686466 397394 686478
rect 432814 686466 433394 686478
rect 468814 686466 469394 686478
rect 504814 686466 505394 686478
rect 540814 686466 541394 686478
rect 576814 686466 577394 686478
rect 585330 686466 585910 686478
rect -2906 686454 586830 686466
rect -2906 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586830 686454
rect -2906 686134 586830 686218
rect -2906 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586830 686134
rect -2906 685886 586830 685898
rect -1986 685874 -1406 685886
rect 814 685874 1394 685886
rect 36814 685874 37394 685886
rect 72814 685874 73394 685886
rect 108814 685874 109394 685886
rect 144814 685874 145394 685886
rect 180814 685874 181394 685886
rect 216814 685874 217394 685886
rect 252814 685874 253394 685886
rect 288814 685874 289394 685886
rect 324814 685874 325394 685886
rect 360814 685874 361394 685886
rect 396814 685874 397394 685886
rect 432814 685874 433394 685886
rect 468814 685874 469394 685886
rect 504814 685874 505394 685886
rect 540814 685874 541394 685886
rect 576814 685874 577394 685886
rect 585330 685874 585910 685886
rect -8426 678906 -7846 678918
rect 29254 678906 29834 678918
rect 65254 678906 65834 678918
rect 101254 678906 101834 678918
rect 137254 678906 137834 678918
rect 173254 678906 173834 678918
rect 209254 678906 209834 678918
rect 245254 678906 245834 678918
rect 281254 678906 281834 678918
rect 317254 678906 317834 678918
rect 353254 678906 353834 678918
rect 389254 678906 389834 678918
rect 425254 678906 425834 678918
rect 461254 678906 461834 678918
rect 497254 678906 497834 678918
rect 533254 678906 533834 678918
rect 569254 678906 569834 678918
rect 591770 678906 592350 678918
rect -8426 678894 592350 678906
rect -8426 678658 -8254 678894
rect -8018 678658 29426 678894
rect 29662 678658 65426 678894
rect 65662 678658 101426 678894
rect 101662 678658 137426 678894
rect 137662 678658 173426 678894
rect 173662 678658 209426 678894
rect 209662 678658 245426 678894
rect 245662 678658 281426 678894
rect 281662 678658 317426 678894
rect 317662 678658 353426 678894
rect 353662 678658 389426 678894
rect 389662 678658 425426 678894
rect 425662 678658 461426 678894
rect 461662 678658 497426 678894
rect 497662 678658 533426 678894
rect 533662 678658 569426 678894
rect 569662 678658 591942 678894
rect 592178 678658 592350 678894
rect -8426 678574 592350 678658
rect -8426 678338 -8254 678574
rect -8018 678338 29426 678574
rect 29662 678338 65426 678574
rect 65662 678338 101426 678574
rect 101662 678338 137426 678574
rect 137662 678338 173426 678574
rect 173662 678338 209426 678574
rect 209662 678338 245426 678574
rect 245662 678338 281426 678574
rect 281662 678338 317426 678574
rect 317662 678338 353426 678574
rect 353662 678338 389426 678574
rect 389662 678338 425426 678574
rect 425662 678338 461426 678574
rect 461662 678338 497426 678574
rect 497662 678338 533426 678574
rect 533662 678338 569426 678574
rect 569662 678338 591942 678574
rect 592178 678338 592350 678574
rect -8426 678326 592350 678338
rect -8426 678314 -7846 678326
rect 29254 678314 29834 678326
rect 65254 678314 65834 678326
rect 101254 678314 101834 678326
rect 137254 678314 137834 678326
rect 173254 678314 173834 678326
rect 209254 678314 209834 678326
rect 245254 678314 245834 678326
rect 281254 678314 281834 678326
rect 317254 678314 317834 678326
rect 353254 678314 353834 678326
rect 389254 678314 389834 678326
rect 425254 678314 425834 678326
rect 461254 678314 461834 678326
rect 497254 678314 497834 678326
rect 533254 678314 533834 678326
rect 569254 678314 569834 678326
rect 591770 678314 592350 678326
rect -6586 675426 -6006 675438
rect 25774 675426 26354 675438
rect 61774 675426 62354 675438
rect 97774 675426 98354 675438
rect 133774 675426 134354 675438
rect 169774 675426 170354 675438
rect 205774 675426 206354 675438
rect 241774 675426 242354 675438
rect 277774 675426 278354 675438
rect 313774 675426 314354 675438
rect 349774 675426 350354 675438
rect 385774 675426 386354 675438
rect 421774 675426 422354 675438
rect 457774 675426 458354 675438
rect 493774 675426 494354 675438
rect 529774 675426 530354 675438
rect 565774 675426 566354 675438
rect 589930 675426 590510 675438
rect -6586 675414 590510 675426
rect -6586 675178 -6414 675414
rect -6178 675178 25946 675414
rect 26182 675178 61946 675414
rect 62182 675178 97946 675414
rect 98182 675178 133946 675414
rect 134182 675178 169946 675414
rect 170182 675178 205946 675414
rect 206182 675178 241946 675414
rect 242182 675178 277946 675414
rect 278182 675178 313946 675414
rect 314182 675178 349946 675414
rect 350182 675178 385946 675414
rect 386182 675178 421946 675414
rect 422182 675178 457946 675414
rect 458182 675178 493946 675414
rect 494182 675178 529946 675414
rect 530182 675178 565946 675414
rect 566182 675178 590102 675414
rect 590338 675178 590510 675414
rect -6586 675094 590510 675178
rect -6586 674858 -6414 675094
rect -6178 674858 25946 675094
rect 26182 674858 61946 675094
rect 62182 674858 97946 675094
rect 98182 674858 133946 675094
rect 134182 674858 169946 675094
rect 170182 674858 205946 675094
rect 206182 674858 241946 675094
rect 242182 674858 277946 675094
rect 278182 674858 313946 675094
rect 314182 674858 349946 675094
rect 350182 674858 385946 675094
rect 386182 674858 421946 675094
rect 422182 674858 457946 675094
rect 458182 674858 493946 675094
rect 494182 674858 529946 675094
rect 530182 674858 565946 675094
rect 566182 674858 590102 675094
rect 590338 674858 590510 675094
rect -6586 674846 590510 674858
rect -6586 674834 -6006 674846
rect 25774 674834 26354 674846
rect 61774 674834 62354 674846
rect 97774 674834 98354 674846
rect 133774 674834 134354 674846
rect 169774 674834 170354 674846
rect 205774 674834 206354 674846
rect 241774 674834 242354 674846
rect 277774 674834 278354 674846
rect 313774 674834 314354 674846
rect 349774 674834 350354 674846
rect 385774 674834 386354 674846
rect 421774 674834 422354 674846
rect 457774 674834 458354 674846
rect 493774 674834 494354 674846
rect 529774 674834 530354 674846
rect 565774 674834 566354 674846
rect 589930 674834 590510 674846
rect -4746 671946 -4166 671958
rect 22294 671946 22874 671958
rect 58294 671946 58874 671958
rect 94294 671946 94874 671958
rect 130294 671946 130874 671958
rect 166294 671946 166874 671958
rect 202294 671946 202874 671958
rect 238294 671946 238874 671958
rect 274294 671946 274874 671958
rect 310294 671946 310874 671958
rect 346294 671946 346874 671958
rect 382294 671946 382874 671958
rect 418294 671946 418874 671958
rect 454294 671946 454874 671958
rect 490294 671946 490874 671958
rect 526294 671946 526874 671958
rect 562294 671946 562874 671958
rect 588090 671946 588670 671958
rect -4746 671934 588670 671946
rect -4746 671698 -4574 671934
rect -4338 671698 22466 671934
rect 22702 671698 58466 671934
rect 58702 671698 94466 671934
rect 94702 671698 130466 671934
rect 130702 671698 166466 671934
rect 166702 671698 202466 671934
rect 202702 671698 238466 671934
rect 238702 671698 274466 671934
rect 274702 671698 310466 671934
rect 310702 671698 346466 671934
rect 346702 671698 382466 671934
rect 382702 671698 418466 671934
rect 418702 671698 454466 671934
rect 454702 671698 490466 671934
rect 490702 671698 526466 671934
rect 526702 671698 562466 671934
rect 562702 671698 588262 671934
rect 588498 671698 588670 671934
rect -4746 671614 588670 671698
rect -4746 671378 -4574 671614
rect -4338 671378 22466 671614
rect 22702 671378 58466 671614
rect 58702 671378 94466 671614
rect 94702 671378 130466 671614
rect 130702 671378 166466 671614
rect 166702 671378 202466 671614
rect 202702 671378 238466 671614
rect 238702 671378 274466 671614
rect 274702 671378 310466 671614
rect 310702 671378 346466 671614
rect 346702 671378 382466 671614
rect 382702 671378 418466 671614
rect 418702 671378 454466 671614
rect 454702 671378 490466 671614
rect 490702 671378 526466 671614
rect 526702 671378 562466 671614
rect 562702 671378 588262 671614
rect 588498 671378 588670 671614
rect -4746 671366 588670 671378
rect -4746 671354 -4166 671366
rect 22294 671354 22874 671366
rect 58294 671354 58874 671366
rect 94294 671354 94874 671366
rect 130294 671354 130874 671366
rect 166294 671354 166874 671366
rect 202294 671354 202874 671366
rect 238294 671354 238874 671366
rect 274294 671354 274874 671366
rect 310294 671354 310874 671366
rect 346294 671354 346874 671366
rect 382294 671354 382874 671366
rect 418294 671354 418874 671366
rect 454294 671354 454874 671366
rect 490294 671354 490874 671366
rect 526294 671354 526874 671366
rect 562294 671354 562874 671366
rect 588090 671354 588670 671366
rect -2906 668466 -2326 668478
rect 18814 668466 19394 668478
rect 54814 668466 55394 668478
rect 90814 668466 91394 668478
rect 126814 668466 127394 668478
rect 162814 668466 163394 668478
rect 198814 668466 199394 668478
rect 234814 668466 235394 668478
rect 270814 668466 271394 668478
rect 306814 668466 307394 668478
rect 342814 668466 343394 668478
rect 378814 668466 379394 668478
rect 414814 668466 415394 668478
rect 450814 668466 451394 668478
rect 486814 668466 487394 668478
rect 522814 668466 523394 668478
rect 558814 668466 559394 668478
rect 586250 668466 586830 668478
rect -2906 668454 586830 668466
rect -2906 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586830 668454
rect -2906 668134 586830 668218
rect -2906 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586830 668134
rect -2906 667886 586830 667898
rect -2906 667874 -2326 667886
rect 18814 667874 19394 667886
rect 54814 667874 55394 667886
rect 90814 667874 91394 667886
rect 126814 667874 127394 667886
rect 162814 667874 163394 667886
rect 198814 667874 199394 667886
rect 234814 667874 235394 667886
rect 270814 667874 271394 667886
rect 306814 667874 307394 667886
rect 342814 667874 343394 667886
rect 378814 667874 379394 667886
rect 414814 667874 415394 667886
rect 450814 667874 451394 667886
rect 486814 667874 487394 667886
rect 522814 667874 523394 667886
rect 558814 667874 559394 667886
rect 586250 667874 586830 667886
rect -7506 660906 -6926 660918
rect 11254 660906 11834 660918
rect 47254 660906 47834 660918
rect 83254 660906 83834 660918
rect 119254 660906 119834 660918
rect 155254 660906 155834 660918
rect 191254 660906 191834 660918
rect 227254 660906 227834 660918
rect 263254 660906 263834 660918
rect 299254 660906 299834 660918
rect 335254 660906 335834 660918
rect 371254 660906 371834 660918
rect 407254 660906 407834 660918
rect 443254 660906 443834 660918
rect 479254 660906 479834 660918
rect 515254 660906 515834 660918
rect 551254 660906 551834 660918
rect 590850 660906 591430 660918
rect -8426 660894 592350 660906
rect -8426 660658 -7334 660894
rect -7098 660658 11426 660894
rect 11662 660658 47426 660894
rect 47662 660658 83426 660894
rect 83662 660658 119426 660894
rect 119662 660658 155426 660894
rect 155662 660658 191426 660894
rect 191662 660658 227426 660894
rect 227662 660658 263426 660894
rect 263662 660658 299426 660894
rect 299662 660658 335426 660894
rect 335662 660658 371426 660894
rect 371662 660658 407426 660894
rect 407662 660658 443426 660894
rect 443662 660658 479426 660894
rect 479662 660658 515426 660894
rect 515662 660658 551426 660894
rect 551662 660658 591022 660894
rect 591258 660658 592350 660894
rect -8426 660574 592350 660658
rect -8426 660338 -7334 660574
rect -7098 660338 11426 660574
rect 11662 660338 47426 660574
rect 47662 660338 83426 660574
rect 83662 660338 119426 660574
rect 119662 660338 155426 660574
rect 155662 660338 191426 660574
rect 191662 660338 227426 660574
rect 227662 660338 263426 660574
rect 263662 660338 299426 660574
rect 299662 660338 335426 660574
rect 335662 660338 371426 660574
rect 371662 660338 407426 660574
rect 407662 660338 443426 660574
rect 443662 660338 479426 660574
rect 479662 660338 515426 660574
rect 515662 660338 551426 660574
rect 551662 660338 591022 660574
rect 591258 660338 592350 660574
rect -8426 660326 592350 660338
rect -7506 660314 -6926 660326
rect 11254 660314 11834 660326
rect 47254 660314 47834 660326
rect 83254 660314 83834 660326
rect 119254 660314 119834 660326
rect 155254 660314 155834 660326
rect 191254 660314 191834 660326
rect 227254 660314 227834 660326
rect 263254 660314 263834 660326
rect 299254 660314 299834 660326
rect 335254 660314 335834 660326
rect 371254 660314 371834 660326
rect 407254 660314 407834 660326
rect 443254 660314 443834 660326
rect 479254 660314 479834 660326
rect 515254 660314 515834 660326
rect 551254 660314 551834 660326
rect 590850 660314 591430 660326
rect -5666 657426 -5086 657438
rect 7774 657426 8354 657438
rect 43774 657426 44354 657438
rect 79774 657426 80354 657438
rect 115774 657426 116354 657438
rect 151774 657426 152354 657438
rect 187774 657426 188354 657438
rect 223774 657426 224354 657438
rect 259774 657426 260354 657438
rect 295774 657426 296354 657438
rect 331774 657426 332354 657438
rect 367774 657426 368354 657438
rect 403774 657426 404354 657438
rect 439774 657426 440354 657438
rect 475774 657426 476354 657438
rect 511774 657426 512354 657438
rect 547774 657426 548354 657438
rect 589010 657426 589590 657438
rect -6586 657414 590510 657426
rect -6586 657178 -5494 657414
rect -5258 657178 7946 657414
rect 8182 657178 43946 657414
rect 44182 657178 79946 657414
rect 80182 657178 115946 657414
rect 116182 657178 151946 657414
rect 152182 657178 187946 657414
rect 188182 657178 223946 657414
rect 224182 657178 259946 657414
rect 260182 657178 295946 657414
rect 296182 657178 331946 657414
rect 332182 657178 367946 657414
rect 368182 657178 403946 657414
rect 404182 657178 439946 657414
rect 440182 657178 475946 657414
rect 476182 657178 511946 657414
rect 512182 657178 547946 657414
rect 548182 657178 589182 657414
rect 589418 657178 590510 657414
rect -6586 657094 590510 657178
rect -6586 656858 -5494 657094
rect -5258 656858 7946 657094
rect 8182 656858 43946 657094
rect 44182 656858 79946 657094
rect 80182 656858 115946 657094
rect 116182 656858 151946 657094
rect 152182 656858 187946 657094
rect 188182 656858 223946 657094
rect 224182 656858 259946 657094
rect 260182 656858 295946 657094
rect 296182 656858 331946 657094
rect 332182 656858 367946 657094
rect 368182 656858 403946 657094
rect 404182 656858 439946 657094
rect 440182 656858 475946 657094
rect 476182 656858 511946 657094
rect 512182 656858 547946 657094
rect 548182 656858 589182 657094
rect 589418 656858 590510 657094
rect -6586 656846 590510 656858
rect -5666 656834 -5086 656846
rect 7774 656834 8354 656846
rect 43774 656834 44354 656846
rect 79774 656834 80354 656846
rect 115774 656834 116354 656846
rect 151774 656834 152354 656846
rect 187774 656834 188354 656846
rect 223774 656834 224354 656846
rect 259774 656834 260354 656846
rect 295774 656834 296354 656846
rect 331774 656834 332354 656846
rect 367774 656834 368354 656846
rect 403774 656834 404354 656846
rect 439774 656834 440354 656846
rect 475774 656834 476354 656846
rect 511774 656834 512354 656846
rect 547774 656834 548354 656846
rect 589010 656834 589590 656846
rect -3826 653946 -3246 653958
rect 4294 653946 4874 653958
rect 40294 653946 40874 653958
rect 76294 653946 76874 653958
rect 112294 653946 112874 653958
rect 148294 653946 148874 653958
rect 184294 653946 184874 653958
rect 220294 653946 220874 653958
rect 256294 653946 256874 653958
rect 292294 653946 292874 653958
rect 328294 653946 328874 653958
rect 364294 653946 364874 653958
rect 400294 653946 400874 653958
rect 436294 653946 436874 653958
rect 472294 653946 472874 653958
rect 508294 653946 508874 653958
rect 544294 653946 544874 653958
rect 580294 653946 580874 653958
rect 587170 653946 587750 653958
rect -4746 653934 588670 653946
rect -4746 653698 -3654 653934
rect -3418 653698 4466 653934
rect 4702 653698 40466 653934
rect 40702 653698 76466 653934
rect 76702 653698 112466 653934
rect 112702 653698 148466 653934
rect 148702 653698 184466 653934
rect 184702 653698 220466 653934
rect 220702 653698 256466 653934
rect 256702 653698 292466 653934
rect 292702 653698 328466 653934
rect 328702 653698 364466 653934
rect 364702 653698 400466 653934
rect 400702 653698 436466 653934
rect 436702 653698 472466 653934
rect 472702 653698 508466 653934
rect 508702 653698 544466 653934
rect 544702 653698 580466 653934
rect 580702 653698 587342 653934
rect 587578 653698 588670 653934
rect -4746 653614 588670 653698
rect -4746 653378 -3654 653614
rect -3418 653378 4466 653614
rect 4702 653378 40466 653614
rect 40702 653378 76466 653614
rect 76702 653378 112466 653614
rect 112702 653378 148466 653614
rect 148702 653378 184466 653614
rect 184702 653378 220466 653614
rect 220702 653378 256466 653614
rect 256702 653378 292466 653614
rect 292702 653378 328466 653614
rect 328702 653378 364466 653614
rect 364702 653378 400466 653614
rect 400702 653378 436466 653614
rect 436702 653378 472466 653614
rect 472702 653378 508466 653614
rect 508702 653378 544466 653614
rect 544702 653378 580466 653614
rect 580702 653378 587342 653614
rect 587578 653378 588670 653614
rect -4746 653366 588670 653378
rect -3826 653354 -3246 653366
rect 4294 653354 4874 653366
rect 40294 653354 40874 653366
rect 76294 653354 76874 653366
rect 112294 653354 112874 653366
rect 148294 653354 148874 653366
rect 184294 653354 184874 653366
rect 220294 653354 220874 653366
rect 256294 653354 256874 653366
rect 292294 653354 292874 653366
rect 328294 653354 328874 653366
rect 364294 653354 364874 653366
rect 400294 653354 400874 653366
rect 436294 653354 436874 653366
rect 472294 653354 472874 653366
rect 508294 653354 508874 653366
rect 544294 653354 544874 653366
rect 580294 653354 580874 653366
rect 587170 653354 587750 653366
rect -1986 650466 -1406 650478
rect 814 650466 1394 650478
rect 36814 650466 37394 650478
rect 72814 650466 73394 650478
rect 108814 650466 109394 650478
rect 144814 650466 145394 650478
rect 180814 650466 181394 650478
rect 216814 650466 217394 650478
rect 252814 650466 253394 650478
rect 288814 650466 289394 650478
rect 324814 650466 325394 650478
rect 360814 650466 361394 650478
rect 396814 650466 397394 650478
rect 432814 650466 433394 650478
rect 468814 650466 469394 650478
rect 504814 650466 505394 650478
rect 540814 650466 541394 650478
rect 576814 650466 577394 650478
rect 585330 650466 585910 650478
rect -2906 650454 586830 650466
rect -2906 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586830 650454
rect -2906 650134 586830 650218
rect -2906 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586830 650134
rect -2906 649886 586830 649898
rect -1986 649874 -1406 649886
rect 814 649874 1394 649886
rect 36814 649874 37394 649886
rect 72814 649874 73394 649886
rect 108814 649874 109394 649886
rect 144814 649874 145394 649886
rect 180814 649874 181394 649886
rect 216814 649874 217394 649886
rect 252814 649874 253394 649886
rect 288814 649874 289394 649886
rect 324814 649874 325394 649886
rect 360814 649874 361394 649886
rect 396814 649874 397394 649886
rect 432814 649874 433394 649886
rect 468814 649874 469394 649886
rect 504814 649874 505394 649886
rect 540814 649874 541394 649886
rect 576814 649874 577394 649886
rect 585330 649874 585910 649886
rect -8426 642906 -7846 642918
rect 29254 642906 29834 642918
rect 65254 642906 65834 642918
rect 101254 642906 101834 642918
rect 137254 642906 137834 642918
rect 173254 642906 173834 642918
rect 209254 642906 209834 642918
rect 245254 642906 245834 642918
rect 281254 642906 281834 642918
rect 317254 642906 317834 642918
rect 353254 642906 353834 642918
rect 389254 642906 389834 642918
rect 425254 642906 425834 642918
rect 461254 642906 461834 642918
rect 497254 642906 497834 642918
rect 533254 642906 533834 642918
rect 569254 642906 569834 642918
rect 591770 642906 592350 642918
rect -8426 642894 592350 642906
rect -8426 642658 -8254 642894
rect -8018 642658 29426 642894
rect 29662 642658 65426 642894
rect 65662 642658 101426 642894
rect 101662 642658 137426 642894
rect 137662 642658 173426 642894
rect 173662 642658 209426 642894
rect 209662 642658 245426 642894
rect 245662 642658 281426 642894
rect 281662 642658 317426 642894
rect 317662 642658 353426 642894
rect 353662 642658 389426 642894
rect 389662 642658 425426 642894
rect 425662 642658 461426 642894
rect 461662 642658 497426 642894
rect 497662 642658 533426 642894
rect 533662 642658 569426 642894
rect 569662 642658 591942 642894
rect 592178 642658 592350 642894
rect -8426 642574 592350 642658
rect -8426 642338 -8254 642574
rect -8018 642338 29426 642574
rect 29662 642338 65426 642574
rect 65662 642338 101426 642574
rect 101662 642338 137426 642574
rect 137662 642338 173426 642574
rect 173662 642338 209426 642574
rect 209662 642338 245426 642574
rect 245662 642338 281426 642574
rect 281662 642338 317426 642574
rect 317662 642338 353426 642574
rect 353662 642338 389426 642574
rect 389662 642338 425426 642574
rect 425662 642338 461426 642574
rect 461662 642338 497426 642574
rect 497662 642338 533426 642574
rect 533662 642338 569426 642574
rect 569662 642338 591942 642574
rect 592178 642338 592350 642574
rect -8426 642326 592350 642338
rect -8426 642314 -7846 642326
rect 29254 642314 29834 642326
rect 65254 642314 65834 642326
rect 101254 642314 101834 642326
rect 137254 642314 137834 642326
rect 173254 642314 173834 642326
rect 209254 642314 209834 642326
rect 245254 642314 245834 642326
rect 281254 642314 281834 642326
rect 317254 642314 317834 642326
rect 353254 642314 353834 642326
rect 389254 642314 389834 642326
rect 425254 642314 425834 642326
rect 461254 642314 461834 642326
rect 497254 642314 497834 642326
rect 533254 642314 533834 642326
rect 569254 642314 569834 642326
rect 591770 642314 592350 642326
rect -6586 639426 -6006 639438
rect 25774 639426 26354 639438
rect 61774 639426 62354 639438
rect 97774 639426 98354 639438
rect 133774 639426 134354 639438
rect 169774 639426 170354 639438
rect 205774 639426 206354 639438
rect 241774 639426 242354 639438
rect 277774 639426 278354 639438
rect 313774 639426 314354 639438
rect 349774 639426 350354 639438
rect 385774 639426 386354 639438
rect 421774 639426 422354 639438
rect 457774 639426 458354 639438
rect 493774 639426 494354 639438
rect 529774 639426 530354 639438
rect 565774 639426 566354 639438
rect 589930 639426 590510 639438
rect -6586 639414 590510 639426
rect -6586 639178 -6414 639414
rect -6178 639178 25946 639414
rect 26182 639178 61946 639414
rect 62182 639178 97946 639414
rect 98182 639178 133946 639414
rect 134182 639178 169946 639414
rect 170182 639178 205946 639414
rect 206182 639178 241946 639414
rect 242182 639178 277946 639414
rect 278182 639178 313946 639414
rect 314182 639178 349946 639414
rect 350182 639178 385946 639414
rect 386182 639178 421946 639414
rect 422182 639178 457946 639414
rect 458182 639178 493946 639414
rect 494182 639178 529946 639414
rect 530182 639178 565946 639414
rect 566182 639178 590102 639414
rect 590338 639178 590510 639414
rect -6586 639094 590510 639178
rect -6586 638858 -6414 639094
rect -6178 638858 25946 639094
rect 26182 638858 61946 639094
rect 62182 638858 97946 639094
rect 98182 638858 133946 639094
rect 134182 638858 169946 639094
rect 170182 638858 205946 639094
rect 206182 638858 241946 639094
rect 242182 638858 277946 639094
rect 278182 638858 313946 639094
rect 314182 638858 349946 639094
rect 350182 638858 385946 639094
rect 386182 638858 421946 639094
rect 422182 638858 457946 639094
rect 458182 638858 493946 639094
rect 494182 638858 529946 639094
rect 530182 638858 565946 639094
rect 566182 638858 590102 639094
rect 590338 638858 590510 639094
rect -6586 638846 590510 638858
rect -6586 638834 -6006 638846
rect 25774 638834 26354 638846
rect 61774 638834 62354 638846
rect 97774 638834 98354 638846
rect 133774 638834 134354 638846
rect 169774 638834 170354 638846
rect 205774 638834 206354 638846
rect 241774 638834 242354 638846
rect 277774 638834 278354 638846
rect 313774 638834 314354 638846
rect 349774 638834 350354 638846
rect 385774 638834 386354 638846
rect 421774 638834 422354 638846
rect 457774 638834 458354 638846
rect 493774 638834 494354 638846
rect 529774 638834 530354 638846
rect 565774 638834 566354 638846
rect 589930 638834 590510 638846
rect -4746 635946 -4166 635958
rect 22294 635946 22874 635958
rect 58294 635946 58874 635958
rect 94294 635946 94874 635958
rect 130294 635946 130874 635958
rect 166294 635946 166874 635958
rect 202294 635946 202874 635958
rect 238294 635946 238874 635958
rect 274294 635946 274874 635958
rect 310294 635946 310874 635958
rect 346294 635946 346874 635958
rect 382294 635946 382874 635958
rect 418294 635946 418874 635958
rect 454294 635946 454874 635958
rect 490294 635946 490874 635958
rect 526294 635946 526874 635958
rect 562294 635946 562874 635958
rect 588090 635946 588670 635958
rect -4746 635934 588670 635946
rect -4746 635698 -4574 635934
rect -4338 635698 22466 635934
rect 22702 635698 58466 635934
rect 58702 635698 94466 635934
rect 94702 635698 130466 635934
rect 130702 635698 166466 635934
rect 166702 635698 202466 635934
rect 202702 635698 238466 635934
rect 238702 635698 274466 635934
rect 274702 635698 310466 635934
rect 310702 635698 346466 635934
rect 346702 635698 382466 635934
rect 382702 635698 418466 635934
rect 418702 635698 454466 635934
rect 454702 635698 490466 635934
rect 490702 635698 526466 635934
rect 526702 635698 562466 635934
rect 562702 635698 588262 635934
rect 588498 635698 588670 635934
rect -4746 635614 588670 635698
rect -4746 635378 -4574 635614
rect -4338 635378 22466 635614
rect 22702 635378 58466 635614
rect 58702 635378 94466 635614
rect 94702 635378 130466 635614
rect 130702 635378 166466 635614
rect 166702 635378 202466 635614
rect 202702 635378 238466 635614
rect 238702 635378 274466 635614
rect 274702 635378 310466 635614
rect 310702 635378 346466 635614
rect 346702 635378 382466 635614
rect 382702 635378 418466 635614
rect 418702 635378 454466 635614
rect 454702 635378 490466 635614
rect 490702 635378 526466 635614
rect 526702 635378 562466 635614
rect 562702 635378 588262 635614
rect 588498 635378 588670 635614
rect -4746 635366 588670 635378
rect -4746 635354 -4166 635366
rect 22294 635354 22874 635366
rect 58294 635354 58874 635366
rect 94294 635354 94874 635366
rect 130294 635354 130874 635366
rect 166294 635354 166874 635366
rect 202294 635354 202874 635366
rect 238294 635354 238874 635366
rect 274294 635354 274874 635366
rect 310294 635354 310874 635366
rect 346294 635354 346874 635366
rect 382294 635354 382874 635366
rect 418294 635354 418874 635366
rect 454294 635354 454874 635366
rect 490294 635354 490874 635366
rect 526294 635354 526874 635366
rect 562294 635354 562874 635366
rect 588090 635354 588670 635366
rect -2906 632466 -2326 632478
rect 18814 632466 19394 632478
rect 54814 632466 55394 632478
rect 90814 632466 91394 632478
rect 126814 632466 127394 632478
rect 162814 632466 163394 632478
rect 198814 632466 199394 632478
rect 234814 632466 235394 632478
rect 270814 632466 271394 632478
rect 306814 632466 307394 632478
rect 342814 632466 343394 632478
rect 378814 632466 379394 632478
rect 414814 632466 415394 632478
rect 450814 632466 451394 632478
rect 486814 632466 487394 632478
rect 522814 632466 523394 632478
rect 558814 632466 559394 632478
rect 586250 632466 586830 632478
rect -2906 632454 586830 632466
rect -2906 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586830 632454
rect -2906 632134 586830 632218
rect -2906 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586830 632134
rect -2906 631886 586830 631898
rect -2906 631874 -2326 631886
rect 18814 631874 19394 631886
rect 54814 631874 55394 631886
rect 90814 631874 91394 631886
rect 126814 631874 127394 631886
rect 162814 631874 163394 631886
rect 198814 631874 199394 631886
rect 234814 631874 235394 631886
rect 270814 631874 271394 631886
rect 306814 631874 307394 631886
rect 342814 631874 343394 631886
rect 378814 631874 379394 631886
rect 414814 631874 415394 631886
rect 450814 631874 451394 631886
rect 486814 631874 487394 631886
rect 522814 631874 523394 631886
rect 558814 631874 559394 631886
rect 586250 631874 586830 631886
rect -7506 624906 -6926 624918
rect 11254 624906 11834 624918
rect 47254 624906 47834 624918
rect 83254 624906 83834 624918
rect 119254 624906 119834 624918
rect 155254 624906 155834 624918
rect 191254 624906 191834 624918
rect 227254 624906 227834 624918
rect 263254 624906 263834 624918
rect 299254 624906 299834 624918
rect 335254 624906 335834 624918
rect 371254 624906 371834 624918
rect 407254 624906 407834 624918
rect 443254 624906 443834 624918
rect 479254 624906 479834 624918
rect 515254 624906 515834 624918
rect 551254 624906 551834 624918
rect 590850 624906 591430 624918
rect -8426 624894 592350 624906
rect -8426 624658 -7334 624894
rect -7098 624658 11426 624894
rect 11662 624658 47426 624894
rect 47662 624658 83426 624894
rect 83662 624658 119426 624894
rect 119662 624658 155426 624894
rect 155662 624658 191426 624894
rect 191662 624658 227426 624894
rect 227662 624658 263426 624894
rect 263662 624658 299426 624894
rect 299662 624658 335426 624894
rect 335662 624658 371426 624894
rect 371662 624658 407426 624894
rect 407662 624658 443426 624894
rect 443662 624658 479426 624894
rect 479662 624658 515426 624894
rect 515662 624658 551426 624894
rect 551662 624658 591022 624894
rect 591258 624658 592350 624894
rect -8426 624574 592350 624658
rect -8426 624338 -7334 624574
rect -7098 624338 11426 624574
rect 11662 624338 47426 624574
rect 47662 624338 83426 624574
rect 83662 624338 119426 624574
rect 119662 624338 155426 624574
rect 155662 624338 191426 624574
rect 191662 624338 227426 624574
rect 227662 624338 263426 624574
rect 263662 624338 299426 624574
rect 299662 624338 335426 624574
rect 335662 624338 371426 624574
rect 371662 624338 407426 624574
rect 407662 624338 443426 624574
rect 443662 624338 479426 624574
rect 479662 624338 515426 624574
rect 515662 624338 551426 624574
rect 551662 624338 591022 624574
rect 591258 624338 592350 624574
rect -8426 624326 592350 624338
rect -7506 624314 -6926 624326
rect 11254 624314 11834 624326
rect 47254 624314 47834 624326
rect 83254 624314 83834 624326
rect 119254 624314 119834 624326
rect 155254 624314 155834 624326
rect 191254 624314 191834 624326
rect 227254 624314 227834 624326
rect 263254 624314 263834 624326
rect 299254 624314 299834 624326
rect 335254 624314 335834 624326
rect 371254 624314 371834 624326
rect 407254 624314 407834 624326
rect 443254 624314 443834 624326
rect 479254 624314 479834 624326
rect 515254 624314 515834 624326
rect 551254 624314 551834 624326
rect 590850 624314 591430 624326
rect -5666 621426 -5086 621438
rect 7774 621426 8354 621438
rect 43774 621426 44354 621438
rect 79774 621426 80354 621438
rect 115774 621426 116354 621438
rect 151774 621426 152354 621438
rect 187774 621426 188354 621438
rect 223774 621426 224354 621438
rect 259774 621426 260354 621438
rect 295774 621426 296354 621438
rect 331774 621426 332354 621438
rect 367774 621426 368354 621438
rect 403774 621426 404354 621438
rect 439774 621426 440354 621438
rect 475774 621426 476354 621438
rect 511774 621426 512354 621438
rect 547774 621426 548354 621438
rect 589010 621426 589590 621438
rect -6586 621414 590510 621426
rect -6586 621178 -5494 621414
rect -5258 621178 7946 621414
rect 8182 621178 43946 621414
rect 44182 621178 79946 621414
rect 80182 621178 115946 621414
rect 116182 621178 151946 621414
rect 152182 621178 187946 621414
rect 188182 621178 223946 621414
rect 224182 621178 259946 621414
rect 260182 621178 295946 621414
rect 296182 621178 331946 621414
rect 332182 621178 367946 621414
rect 368182 621178 403946 621414
rect 404182 621178 439946 621414
rect 440182 621178 475946 621414
rect 476182 621178 511946 621414
rect 512182 621178 547946 621414
rect 548182 621178 589182 621414
rect 589418 621178 590510 621414
rect -6586 621094 590510 621178
rect -6586 620858 -5494 621094
rect -5258 620858 7946 621094
rect 8182 620858 43946 621094
rect 44182 620858 79946 621094
rect 80182 620858 115946 621094
rect 116182 620858 151946 621094
rect 152182 620858 187946 621094
rect 188182 620858 223946 621094
rect 224182 620858 259946 621094
rect 260182 620858 295946 621094
rect 296182 620858 331946 621094
rect 332182 620858 367946 621094
rect 368182 620858 403946 621094
rect 404182 620858 439946 621094
rect 440182 620858 475946 621094
rect 476182 620858 511946 621094
rect 512182 620858 547946 621094
rect 548182 620858 589182 621094
rect 589418 620858 590510 621094
rect -6586 620846 590510 620858
rect -5666 620834 -5086 620846
rect 7774 620834 8354 620846
rect 43774 620834 44354 620846
rect 79774 620834 80354 620846
rect 115774 620834 116354 620846
rect 151774 620834 152354 620846
rect 187774 620834 188354 620846
rect 223774 620834 224354 620846
rect 259774 620834 260354 620846
rect 295774 620834 296354 620846
rect 331774 620834 332354 620846
rect 367774 620834 368354 620846
rect 403774 620834 404354 620846
rect 439774 620834 440354 620846
rect 475774 620834 476354 620846
rect 511774 620834 512354 620846
rect 547774 620834 548354 620846
rect 589010 620834 589590 620846
rect -3826 617946 -3246 617958
rect 4294 617946 4874 617958
rect 40294 617946 40874 617958
rect 76294 617946 76874 617958
rect 112294 617946 112874 617958
rect 148294 617946 148874 617958
rect 184294 617946 184874 617958
rect 220294 617946 220874 617958
rect 256294 617946 256874 617958
rect 292294 617946 292874 617958
rect 328294 617946 328874 617958
rect 364294 617946 364874 617958
rect 400294 617946 400874 617958
rect 436294 617946 436874 617958
rect 472294 617946 472874 617958
rect 508294 617946 508874 617958
rect 544294 617946 544874 617958
rect 580294 617946 580874 617958
rect 587170 617946 587750 617958
rect -4746 617934 588670 617946
rect -4746 617698 -3654 617934
rect -3418 617698 4466 617934
rect 4702 617698 40466 617934
rect 40702 617698 76466 617934
rect 76702 617698 112466 617934
rect 112702 617698 148466 617934
rect 148702 617698 184466 617934
rect 184702 617698 220466 617934
rect 220702 617698 256466 617934
rect 256702 617698 292466 617934
rect 292702 617698 328466 617934
rect 328702 617698 364466 617934
rect 364702 617698 400466 617934
rect 400702 617698 436466 617934
rect 436702 617698 472466 617934
rect 472702 617698 508466 617934
rect 508702 617698 544466 617934
rect 544702 617698 580466 617934
rect 580702 617698 587342 617934
rect 587578 617698 588670 617934
rect -4746 617614 588670 617698
rect -4746 617378 -3654 617614
rect -3418 617378 4466 617614
rect 4702 617378 40466 617614
rect 40702 617378 76466 617614
rect 76702 617378 112466 617614
rect 112702 617378 148466 617614
rect 148702 617378 184466 617614
rect 184702 617378 220466 617614
rect 220702 617378 256466 617614
rect 256702 617378 292466 617614
rect 292702 617378 328466 617614
rect 328702 617378 364466 617614
rect 364702 617378 400466 617614
rect 400702 617378 436466 617614
rect 436702 617378 472466 617614
rect 472702 617378 508466 617614
rect 508702 617378 544466 617614
rect 544702 617378 580466 617614
rect 580702 617378 587342 617614
rect 587578 617378 588670 617614
rect -4746 617366 588670 617378
rect -3826 617354 -3246 617366
rect 4294 617354 4874 617366
rect 40294 617354 40874 617366
rect 76294 617354 76874 617366
rect 112294 617354 112874 617366
rect 148294 617354 148874 617366
rect 184294 617354 184874 617366
rect 220294 617354 220874 617366
rect 256294 617354 256874 617366
rect 292294 617354 292874 617366
rect 328294 617354 328874 617366
rect 364294 617354 364874 617366
rect 400294 617354 400874 617366
rect 436294 617354 436874 617366
rect 472294 617354 472874 617366
rect 508294 617354 508874 617366
rect 544294 617354 544874 617366
rect 580294 617354 580874 617366
rect 587170 617354 587750 617366
rect -1986 614466 -1406 614478
rect 814 614466 1394 614478
rect 36814 614466 37394 614478
rect 72814 614466 73394 614478
rect 108814 614466 109394 614478
rect 144814 614466 145394 614478
rect 180814 614466 181394 614478
rect 216814 614466 217394 614478
rect 252814 614466 253394 614478
rect 288814 614466 289394 614478
rect 324814 614466 325394 614478
rect 360814 614466 361394 614478
rect 396814 614466 397394 614478
rect 432814 614466 433394 614478
rect 468814 614466 469394 614478
rect 504814 614466 505394 614478
rect 540814 614466 541394 614478
rect 576814 614466 577394 614478
rect 585330 614466 585910 614478
rect -2906 614454 586830 614466
rect -2906 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586830 614454
rect -2906 614134 586830 614218
rect -2906 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586830 614134
rect -2906 613886 586830 613898
rect -1986 613874 -1406 613886
rect 814 613874 1394 613886
rect 36814 613874 37394 613886
rect 72814 613874 73394 613886
rect 108814 613874 109394 613886
rect 144814 613874 145394 613886
rect 180814 613874 181394 613886
rect 216814 613874 217394 613886
rect 252814 613874 253394 613886
rect 288814 613874 289394 613886
rect 324814 613874 325394 613886
rect 360814 613874 361394 613886
rect 396814 613874 397394 613886
rect 432814 613874 433394 613886
rect 468814 613874 469394 613886
rect 504814 613874 505394 613886
rect 540814 613874 541394 613886
rect 576814 613874 577394 613886
rect 585330 613874 585910 613886
rect -8426 606906 -7846 606918
rect 29254 606906 29834 606918
rect 65254 606906 65834 606918
rect 101254 606906 101834 606918
rect 137254 606906 137834 606918
rect 173254 606906 173834 606918
rect 209254 606906 209834 606918
rect 245254 606906 245834 606918
rect 281254 606906 281834 606918
rect 317254 606906 317834 606918
rect 353254 606906 353834 606918
rect 389254 606906 389834 606918
rect 425254 606906 425834 606918
rect 461254 606906 461834 606918
rect 497254 606906 497834 606918
rect 533254 606906 533834 606918
rect 569254 606906 569834 606918
rect 591770 606906 592350 606918
rect -8426 606894 592350 606906
rect -8426 606658 -8254 606894
rect -8018 606658 29426 606894
rect 29662 606658 65426 606894
rect 65662 606658 101426 606894
rect 101662 606658 137426 606894
rect 137662 606658 173426 606894
rect 173662 606658 209426 606894
rect 209662 606658 245426 606894
rect 245662 606658 281426 606894
rect 281662 606658 317426 606894
rect 317662 606658 353426 606894
rect 353662 606658 389426 606894
rect 389662 606658 425426 606894
rect 425662 606658 461426 606894
rect 461662 606658 497426 606894
rect 497662 606658 533426 606894
rect 533662 606658 569426 606894
rect 569662 606658 591942 606894
rect 592178 606658 592350 606894
rect -8426 606574 592350 606658
rect -8426 606338 -8254 606574
rect -8018 606338 29426 606574
rect 29662 606338 65426 606574
rect 65662 606338 101426 606574
rect 101662 606338 137426 606574
rect 137662 606338 173426 606574
rect 173662 606338 209426 606574
rect 209662 606338 245426 606574
rect 245662 606338 281426 606574
rect 281662 606338 317426 606574
rect 317662 606338 353426 606574
rect 353662 606338 389426 606574
rect 389662 606338 425426 606574
rect 425662 606338 461426 606574
rect 461662 606338 497426 606574
rect 497662 606338 533426 606574
rect 533662 606338 569426 606574
rect 569662 606338 591942 606574
rect 592178 606338 592350 606574
rect -8426 606326 592350 606338
rect -8426 606314 -7846 606326
rect 29254 606314 29834 606326
rect 65254 606314 65834 606326
rect 101254 606314 101834 606326
rect 137254 606314 137834 606326
rect 173254 606314 173834 606326
rect 209254 606314 209834 606326
rect 245254 606314 245834 606326
rect 281254 606314 281834 606326
rect 317254 606314 317834 606326
rect 353254 606314 353834 606326
rect 389254 606314 389834 606326
rect 425254 606314 425834 606326
rect 461254 606314 461834 606326
rect 497254 606314 497834 606326
rect 533254 606314 533834 606326
rect 569254 606314 569834 606326
rect 591770 606314 592350 606326
rect -6586 603426 -6006 603438
rect 25774 603426 26354 603438
rect 61774 603426 62354 603438
rect 97774 603426 98354 603438
rect 133774 603426 134354 603438
rect 169774 603426 170354 603438
rect 205774 603426 206354 603438
rect 241774 603426 242354 603438
rect 277774 603426 278354 603438
rect 313774 603426 314354 603438
rect 349774 603426 350354 603438
rect 385774 603426 386354 603438
rect 421774 603426 422354 603438
rect 457774 603426 458354 603438
rect 493774 603426 494354 603438
rect 529774 603426 530354 603438
rect 565774 603426 566354 603438
rect 589930 603426 590510 603438
rect -6586 603414 590510 603426
rect -6586 603178 -6414 603414
rect -6178 603178 25946 603414
rect 26182 603178 61946 603414
rect 62182 603178 97946 603414
rect 98182 603178 133946 603414
rect 134182 603178 169946 603414
rect 170182 603178 205946 603414
rect 206182 603178 241946 603414
rect 242182 603178 277946 603414
rect 278182 603178 313946 603414
rect 314182 603178 349946 603414
rect 350182 603178 385946 603414
rect 386182 603178 421946 603414
rect 422182 603178 457946 603414
rect 458182 603178 493946 603414
rect 494182 603178 529946 603414
rect 530182 603178 565946 603414
rect 566182 603178 590102 603414
rect 590338 603178 590510 603414
rect -6586 603094 590510 603178
rect -6586 602858 -6414 603094
rect -6178 602858 25946 603094
rect 26182 602858 61946 603094
rect 62182 602858 97946 603094
rect 98182 602858 133946 603094
rect 134182 602858 169946 603094
rect 170182 602858 205946 603094
rect 206182 602858 241946 603094
rect 242182 602858 277946 603094
rect 278182 602858 313946 603094
rect 314182 602858 349946 603094
rect 350182 602858 385946 603094
rect 386182 602858 421946 603094
rect 422182 602858 457946 603094
rect 458182 602858 493946 603094
rect 494182 602858 529946 603094
rect 530182 602858 565946 603094
rect 566182 602858 590102 603094
rect 590338 602858 590510 603094
rect -6586 602846 590510 602858
rect -6586 602834 -6006 602846
rect 25774 602834 26354 602846
rect 61774 602834 62354 602846
rect 97774 602834 98354 602846
rect 133774 602834 134354 602846
rect 169774 602834 170354 602846
rect 205774 602834 206354 602846
rect 241774 602834 242354 602846
rect 277774 602834 278354 602846
rect 313774 602834 314354 602846
rect 349774 602834 350354 602846
rect 385774 602834 386354 602846
rect 421774 602834 422354 602846
rect 457774 602834 458354 602846
rect 493774 602834 494354 602846
rect 529774 602834 530354 602846
rect 565774 602834 566354 602846
rect 589930 602834 590510 602846
rect -4746 599946 -4166 599958
rect 22294 599946 22874 599958
rect 58294 599946 58874 599958
rect 94294 599946 94874 599958
rect 130294 599946 130874 599958
rect 166294 599946 166874 599958
rect 202294 599946 202874 599958
rect 238294 599946 238874 599958
rect 274294 599946 274874 599958
rect 310294 599946 310874 599958
rect 346294 599946 346874 599958
rect 382294 599946 382874 599958
rect 418294 599946 418874 599958
rect 454294 599946 454874 599958
rect 490294 599946 490874 599958
rect 526294 599946 526874 599958
rect 562294 599946 562874 599958
rect 588090 599946 588670 599958
rect -4746 599934 588670 599946
rect -4746 599698 -4574 599934
rect -4338 599698 22466 599934
rect 22702 599698 58466 599934
rect 58702 599698 94466 599934
rect 94702 599698 130466 599934
rect 130702 599698 166466 599934
rect 166702 599698 202466 599934
rect 202702 599698 238466 599934
rect 238702 599698 274466 599934
rect 274702 599698 310466 599934
rect 310702 599698 346466 599934
rect 346702 599698 382466 599934
rect 382702 599698 418466 599934
rect 418702 599698 454466 599934
rect 454702 599698 490466 599934
rect 490702 599698 526466 599934
rect 526702 599698 562466 599934
rect 562702 599698 588262 599934
rect 588498 599698 588670 599934
rect -4746 599614 588670 599698
rect -4746 599378 -4574 599614
rect -4338 599378 22466 599614
rect 22702 599378 58466 599614
rect 58702 599378 94466 599614
rect 94702 599378 130466 599614
rect 130702 599378 166466 599614
rect 166702 599378 202466 599614
rect 202702 599378 238466 599614
rect 238702 599378 274466 599614
rect 274702 599378 310466 599614
rect 310702 599378 346466 599614
rect 346702 599378 382466 599614
rect 382702 599378 418466 599614
rect 418702 599378 454466 599614
rect 454702 599378 490466 599614
rect 490702 599378 526466 599614
rect 526702 599378 562466 599614
rect 562702 599378 588262 599614
rect 588498 599378 588670 599614
rect -4746 599366 588670 599378
rect -4746 599354 -4166 599366
rect 22294 599354 22874 599366
rect 58294 599354 58874 599366
rect 94294 599354 94874 599366
rect 130294 599354 130874 599366
rect 166294 599354 166874 599366
rect 202294 599354 202874 599366
rect 238294 599354 238874 599366
rect 274294 599354 274874 599366
rect 310294 599354 310874 599366
rect 346294 599354 346874 599366
rect 382294 599354 382874 599366
rect 418294 599354 418874 599366
rect 454294 599354 454874 599366
rect 490294 599354 490874 599366
rect 526294 599354 526874 599366
rect 562294 599354 562874 599366
rect 588090 599354 588670 599366
rect -2906 596466 -2326 596478
rect 18814 596466 19394 596478
rect 54814 596466 55394 596478
rect 90814 596466 91394 596478
rect 126814 596466 127394 596478
rect 162814 596466 163394 596478
rect 198814 596466 199394 596478
rect 234814 596466 235394 596478
rect 270814 596466 271394 596478
rect 306814 596466 307394 596478
rect 342814 596466 343394 596478
rect 378814 596466 379394 596478
rect 414814 596466 415394 596478
rect 450814 596466 451394 596478
rect 486814 596466 487394 596478
rect 522814 596466 523394 596478
rect 558814 596466 559394 596478
rect 586250 596466 586830 596478
rect -2906 596454 586830 596466
rect -2906 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586830 596454
rect -2906 596134 586830 596218
rect -2906 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586830 596134
rect -2906 595886 586830 595898
rect -2906 595874 -2326 595886
rect 18814 595874 19394 595886
rect 54814 595874 55394 595886
rect 90814 595874 91394 595886
rect 126814 595874 127394 595886
rect 162814 595874 163394 595886
rect 198814 595874 199394 595886
rect 234814 595874 235394 595886
rect 270814 595874 271394 595886
rect 306814 595874 307394 595886
rect 342814 595874 343394 595886
rect 378814 595874 379394 595886
rect 414814 595874 415394 595886
rect 450814 595874 451394 595886
rect 486814 595874 487394 595886
rect 522814 595874 523394 595886
rect 558814 595874 559394 595886
rect 586250 595874 586830 595886
rect -7506 588906 -6926 588918
rect 11254 588906 11834 588918
rect 47254 588906 47834 588918
rect 83254 588906 83834 588918
rect 119254 588906 119834 588918
rect 155254 588906 155834 588918
rect 191254 588906 191834 588918
rect 227254 588906 227834 588918
rect 263254 588906 263834 588918
rect 299254 588906 299834 588918
rect 335254 588906 335834 588918
rect 371254 588906 371834 588918
rect 407254 588906 407834 588918
rect 443254 588906 443834 588918
rect 479254 588906 479834 588918
rect 515254 588906 515834 588918
rect 551254 588906 551834 588918
rect 590850 588906 591430 588918
rect -8426 588894 592350 588906
rect -8426 588658 -7334 588894
rect -7098 588658 11426 588894
rect 11662 588658 47426 588894
rect 47662 588658 83426 588894
rect 83662 588658 119426 588894
rect 119662 588658 155426 588894
rect 155662 588658 191426 588894
rect 191662 588658 227426 588894
rect 227662 588658 263426 588894
rect 263662 588658 299426 588894
rect 299662 588658 335426 588894
rect 335662 588658 371426 588894
rect 371662 588658 407426 588894
rect 407662 588658 443426 588894
rect 443662 588658 479426 588894
rect 479662 588658 515426 588894
rect 515662 588658 551426 588894
rect 551662 588658 591022 588894
rect 591258 588658 592350 588894
rect -8426 588574 592350 588658
rect -8426 588338 -7334 588574
rect -7098 588338 11426 588574
rect 11662 588338 47426 588574
rect 47662 588338 83426 588574
rect 83662 588338 119426 588574
rect 119662 588338 155426 588574
rect 155662 588338 191426 588574
rect 191662 588338 227426 588574
rect 227662 588338 263426 588574
rect 263662 588338 299426 588574
rect 299662 588338 335426 588574
rect 335662 588338 371426 588574
rect 371662 588338 407426 588574
rect 407662 588338 443426 588574
rect 443662 588338 479426 588574
rect 479662 588338 515426 588574
rect 515662 588338 551426 588574
rect 551662 588338 591022 588574
rect 591258 588338 592350 588574
rect -8426 588326 592350 588338
rect -7506 588314 -6926 588326
rect 11254 588314 11834 588326
rect 47254 588314 47834 588326
rect 83254 588314 83834 588326
rect 119254 588314 119834 588326
rect 155254 588314 155834 588326
rect 191254 588314 191834 588326
rect 227254 588314 227834 588326
rect 263254 588314 263834 588326
rect 299254 588314 299834 588326
rect 335254 588314 335834 588326
rect 371254 588314 371834 588326
rect 407254 588314 407834 588326
rect 443254 588314 443834 588326
rect 479254 588314 479834 588326
rect 515254 588314 515834 588326
rect 551254 588314 551834 588326
rect 590850 588314 591430 588326
rect -5666 585426 -5086 585438
rect 7774 585426 8354 585438
rect 43774 585426 44354 585438
rect 79774 585426 80354 585438
rect 115774 585426 116354 585438
rect 151774 585426 152354 585438
rect 187774 585426 188354 585438
rect 223774 585426 224354 585438
rect 259774 585426 260354 585438
rect 295774 585426 296354 585438
rect 331774 585426 332354 585438
rect 367774 585426 368354 585438
rect 403774 585426 404354 585438
rect 439774 585426 440354 585438
rect 475774 585426 476354 585438
rect 511774 585426 512354 585438
rect 547774 585426 548354 585438
rect 589010 585426 589590 585438
rect -6586 585414 590510 585426
rect -6586 585178 -5494 585414
rect -5258 585178 7946 585414
rect 8182 585178 43946 585414
rect 44182 585178 79946 585414
rect 80182 585178 115946 585414
rect 116182 585178 151946 585414
rect 152182 585178 187946 585414
rect 188182 585178 223946 585414
rect 224182 585178 259946 585414
rect 260182 585178 295946 585414
rect 296182 585178 331946 585414
rect 332182 585178 367946 585414
rect 368182 585178 403946 585414
rect 404182 585178 439946 585414
rect 440182 585178 475946 585414
rect 476182 585178 511946 585414
rect 512182 585178 547946 585414
rect 548182 585178 589182 585414
rect 589418 585178 590510 585414
rect -6586 585094 590510 585178
rect -6586 584858 -5494 585094
rect -5258 584858 7946 585094
rect 8182 584858 43946 585094
rect 44182 584858 79946 585094
rect 80182 584858 115946 585094
rect 116182 584858 151946 585094
rect 152182 584858 187946 585094
rect 188182 584858 223946 585094
rect 224182 584858 259946 585094
rect 260182 584858 295946 585094
rect 296182 584858 331946 585094
rect 332182 584858 367946 585094
rect 368182 584858 403946 585094
rect 404182 584858 439946 585094
rect 440182 584858 475946 585094
rect 476182 584858 511946 585094
rect 512182 584858 547946 585094
rect 548182 584858 589182 585094
rect 589418 584858 590510 585094
rect -6586 584846 590510 584858
rect -5666 584834 -5086 584846
rect 7774 584834 8354 584846
rect 43774 584834 44354 584846
rect 79774 584834 80354 584846
rect 115774 584834 116354 584846
rect 151774 584834 152354 584846
rect 187774 584834 188354 584846
rect 223774 584834 224354 584846
rect 259774 584834 260354 584846
rect 295774 584834 296354 584846
rect 331774 584834 332354 584846
rect 367774 584834 368354 584846
rect 403774 584834 404354 584846
rect 439774 584834 440354 584846
rect 475774 584834 476354 584846
rect 511774 584834 512354 584846
rect 547774 584834 548354 584846
rect 589010 584834 589590 584846
rect -3826 581946 -3246 581958
rect 4294 581946 4874 581958
rect 40294 581946 40874 581958
rect 76294 581946 76874 581958
rect 112294 581946 112874 581958
rect 148294 581946 148874 581958
rect 184294 581946 184874 581958
rect 220294 581946 220874 581958
rect 256294 581946 256874 581958
rect 292294 581946 292874 581958
rect 328294 581946 328874 581958
rect 364294 581946 364874 581958
rect 400294 581946 400874 581958
rect 436294 581946 436874 581958
rect 472294 581946 472874 581958
rect 508294 581946 508874 581958
rect 544294 581946 544874 581958
rect 580294 581946 580874 581958
rect 587170 581946 587750 581958
rect -4746 581934 588670 581946
rect -4746 581698 -3654 581934
rect -3418 581698 4466 581934
rect 4702 581698 40466 581934
rect 40702 581698 76466 581934
rect 76702 581698 112466 581934
rect 112702 581698 148466 581934
rect 148702 581698 184466 581934
rect 184702 581698 220466 581934
rect 220702 581698 256466 581934
rect 256702 581698 292466 581934
rect 292702 581698 328466 581934
rect 328702 581698 364466 581934
rect 364702 581698 400466 581934
rect 400702 581698 436466 581934
rect 436702 581698 472466 581934
rect 472702 581698 508466 581934
rect 508702 581698 544466 581934
rect 544702 581698 580466 581934
rect 580702 581698 587342 581934
rect 587578 581698 588670 581934
rect -4746 581614 588670 581698
rect -4746 581378 -3654 581614
rect -3418 581378 4466 581614
rect 4702 581378 40466 581614
rect 40702 581378 76466 581614
rect 76702 581378 112466 581614
rect 112702 581378 148466 581614
rect 148702 581378 184466 581614
rect 184702 581378 220466 581614
rect 220702 581378 256466 581614
rect 256702 581378 292466 581614
rect 292702 581378 328466 581614
rect 328702 581378 364466 581614
rect 364702 581378 400466 581614
rect 400702 581378 436466 581614
rect 436702 581378 472466 581614
rect 472702 581378 508466 581614
rect 508702 581378 544466 581614
rect 544702 581378 580466 581614
rect 580702 581378 587342 581614
rect 587578 581378 588670 581614
rect -4746 581366 588670 581378
rect -3826 581354 -3246 581366
rect 4294 581354 4874 581366
rect 40294 581354 40874 581366
rect 76294 581354 76874 581366
rect 112294 581354 112874 581366
rect 148294 581354 148874 581366
rect 184294 581354 184874 581366
rect 220294 581354 220874 581366
rect 256294 581354 256874 581366
rect 292294 581354 292874 581366
rect 328294 581354 328874 581366
rect 364294 581354 364874 581366
rect 400294 581354 400874 581366
rect 436294 581354 436874 581366
rect 472294 581354 472874 581366
rect 508294 581354 508874 581366
rect 544294 581354 544874 581366
rect 580294 581354 580874 581366
rect 587170 581354 587750 581366
rect -1986 578466 -1406 578478
rect 814 578466 1394 578478
rect 36814 578466 37394 578478
rect 72814 578466 73394 578478
rect 108814 578466 109394 578478
rect 144814 578466 145394 578478
rect 180814 578466 181394 578478
rect 216814 578466 217394 578478
rect 252814 578466 253394 578478
rect 288814 578466 289394 578478
rect 324814 578466 325394 578478
rect 360814 578466 361394 578478
rect 396814 578466 397394 578478
rect 432814 578466 433394 578478
rect 468814 578466 469394 578478
rect 504814 578466 505394 578478
rect 540814 578466 541394 578478
rect 576814 578466 577394 578478
rect 585330 578466 585910 578478
rect -2906 578454 586830 578466
rect -2906 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586830 578454
rect -2906 578134 586830 578218
rect -2906 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586830 578134
rect -2906 577886 586830 577898
rect -1986 577874 -1406 577886
rect 814 577874 1394 577886
rect 36814 577874 37394 577886
rect 72814 577874 73394 577886
rect 108814 577874 109394 577886
rect 144814 577874 145394 577886
rect 180814 577874 181394 577886
rect 216814 577874 217394 577886
rect 252814 577874 253394 577886
rect 288814 577874 289394 577886
rect 324814 577874 325394 577886
rect 360814 577874 361394 577886
rect 396814 577874 397394 577886
rect 432814 577874 433394 577886
rect 468814 577874 469394 577886
rect 504814 577874 505394 577886
rect 540814 577874 541394 577886
rect 576814 577874 577394 577886
rect 585330 577874 585910 577886
rect -8426 570906 -7846 570918
rect 29254 570906 29834 570918
rect 65254 570906 65834 570918
rect 101254 570906 101834 570918
rect 137254 570906 137834 570918
rect 173254 570906 173834 570918
rect 209254 570906 209834 570918
rect 245254 570906 245834 570918
rect 281254 570906 281834 570918
rect 317254 570906 317834 570918
rect 353254 570906 353834 570918
rect 389254 570906 389834 570918
rect 425254 570906 425834 570918
rect 461254 570906 461834 570918
rect 497254 570906 497834 570918
rect 533254 570906 533834 570918
rect 569254 570906 569834 570918
rect 591770 570906 592350 570918
rect -8426 570894 592350 570906
rect -8426 570658 -8254 570894
rect -8018 570658 29426 570894
rect 29662 570658 65426 570894
rect 65662 570658 101426 570894
rect 101662 570658 137426 570894
rect 137662 570658 173426 570894
rect 173662 570658 209426 570894
rect 209662 570658 245426 570894
rect 245662 570658 281426 570894
rect 281662 570658 317426 570894
rect 317662 570658 353426 570894
rect 353662 570658 389426 570894
rect 389662 570658 425426 570894
rect 425662 570658 461426 570894
rect 461662 570658 497426 570894
rect 497662 570658 533426 570894
rect 533662 570658 569426 570894
rect 569662 570658 591942 570894
rect 592178 570658 592350 570894
rect -8426 570574 592350 570658
rect -8426 570338 -8254 570574
rect -8018 570338 29426 570574
rect 29662 570338 65426 570574
rect 65662 570338 101426 570574
rect 101662 570338 137426 570574
rect 137662 570338 173426 570574
rect 173662 570338 209426 570574
rect 209662 570338 245426 570574
rect 245662 570338 281426 570574
rect 281662 570338 317426 570574
rect 317662 570338 353426 570574
rect 353662 570338 389426 570574
rect 389662 570338 425426 570574
rect 425662 570338 461426 570574
rect 461662 570338 497426 570574
rect 497662 570338 533426 570574
rect 533662 570338 569426 570574
rect 569662 570338 591942 570574
rect 592178 570338 592350 570574
rect -8426 570326 592350 570338
rect -8426 570314 -7846 570326
rect 29254 570314 29834 570326
rect 65254 570314 65834 570326
rect 101254 570314 101834 570326
rect 137254 570314 137834 570326
rect 173254 570314 173834 570326
rect 209254 570314 209834 570326
rect 245254 570314 245834 570326
rect 281254 570314 281834 570326
rect 317254 570314 317834 570326
rect 353254 570314 353834 570326
rect 389254 570314 389834 570326
rect 425254 570314 425834 570326
rect 461254 570314 461834 570326
rect 497254 570314 497834 570326
rect 533254 570314 533834 570326
rect 569254 570314 569834 570326
rect 591770 570314 592350 570326
rect -6586 567426 -6006 567438
rect 25774 567426 26354 567438
rect 61774 567426 62354 567438
rect 97774 567426 98354 567438
rect 133774 567426 134354 567438
rect 169774 567426 170354 567438
rect 205774 567426 206354 567438
rect 241774 567426 242354 567438
rect 277774 567426 278354 567438
rect 313774 567426 314354 567438
rect 349774 567426 350354 567438
rect 385774 567426 386354 567438
rect 421774 567426 422354 567438
rect 457774 567426 458354 567438
rect 493774 567426 494354 567438
rect 529774 567426 530354 567438
rect 565774 567426 566354 567438
rect 589930 567426 590510 567438
rect -6586 567414 590510 567426
rect -6586 567178 -6414 567414
rect -6178 567178 25946 567414
rect 26182 567178 61946 567414
rect 62182 567178 97946 567414
rect 98182 567178 133946 567414
rect 134182 567178 169946 567414
rect 170182 567178 205946 567414
rect 206182 567178 241946 567414
rect 242182 567178 277946 567414
rect 278182 567178 313946 567414
rect 314182 567178 349946 567414
rect 350182 567178 385946 567414
rect 386182 567178 421946 567414
rect 422182 567178 457946 567414
rect 458182 567178 493946 567414
rect 494182 567178 529946 567414
rect 530182 567178 565946 567414
rect 566182 567178 590102 567414
rect 590338 567178 590510 567414
rect -6586 567094 590510 567178
rect -6586 566858 -6414 567094
rect -6178 566858 25946 567094
rect 26182 566858 61946 567094
rect 62182 566858 97946 567094
rect 98182 566858 133946 567094
rect 134182 566858 169946 567094
rect 170182 566858 205946 567094
rect 206182 566858 241946 567094
rect 242182 566858 277946 567094
rect 278182 566858 313946 567094
rect 314182 566858 349946 567094
rect 350182 566858 385946 567094
rect 386182 566858 421946 567094
rect 422182 566858 457946 567094
rect 458182 566858 493946 567094
rect 494182 566858 529946 567094
rect 530182 566858 565946 567094
rect 566182 566858 590102 567094
rect 590338 566858 590510 567094
rect -6586 566846 590510 566858
rect -6586 566834 -6006 566846
rect 25774 566834 26354 566846
rect 61774 566834 62354 566846
rect 97774 566834 98354 566846
rect 133774 566834 134354 566846
rect 169774 566834 170354 566846
rect 205774 566834 206354 566846
rect 241774 566834 242354 566846
rect 277774 566834 278354 566846
rect 313774 566834 314354 566846
rect 349774 566834 350354 566846
rect 385774 566834 386354 566846
rect 421774 566834 422354 566846
rect 457774 566834 458354 566846
rect 493774 566834 494354 566846
rect 529774 566834 530354 566846
rect 565774 566834 566354 566846
rect 589930 566834 590510 566846
rect -4746 563946 -4166 563958
rect 22294 563946 22874 563958
rect 58294 563946 58874 563958
rect 94294 563946 94874 563958
rect 130294 563946 130874 563958
rect 166294 563946 166874 563958
rect 202294 563946 202874 563958
rect 238294 563946 238874 563958
rect 274294 563946 274874 563958
rect 310294 563946 310874 563958
rect 346294 563946 346874 563958
rect 382294 563946 382874 563958
rect 418294 563946 418874 563958
rect 454294 563946 454874 563958
rect 490294 563946 490874 563958
rect 526294 563946 526874 563958
rect 562294 563946 562874 563958
rect 588090 563946 588670 563958
rect -4746 563934 588670 563946
rect -4746 563698 -4574 563934
rect -4338 563698 22466 563934
rect 22702 563698 58466 563934
rect 58702 563698 94466 563934
rect 94702 563698 130466 563934
rect 130702 563698 166466 563934
rect 166702 563698 202466 563934
rect 202702 563698 238466 563934
rect 238702 563698 274466 563934
rect 274702 563698 310466 563934
rect 310702 563698 346466 563934
rect 346702 563698 382466 563934
rect 382702 563698 418466 563934
rect 418702 563698 454466 563934
rect 454702 563698 490466 563934
rect 490702 563698 526466 563934
rect 526702 563698 562466 563934
rect 562702 563698 588262 563934
rect 588498 563698 588670 563934
rect -4746 563614 588670 563698
rect -4746 563378 -4574 563614
rect -4338 563378 22466 563614
rect 22702 563378 58466 563614
rect 58702 563378 94466 563614
rect 94702 563378 130466 563614
rect 130702 563378 166466 563614
rect 166702 563378 202466 563614
rect 202702 563378 238466 563614
rect 238702 563378 274466 563614
rect 274702 563378 310466 563614
rect 310702 563378 346466 563614
rect 346702 563378 382466 563614
rect 382702 563378 418466 563614
rect 418702 563378 454466 563614
rect 454702 563378 490466 563614
rect 490702 563378 526466 563614
rect 526702 563378 562466 563614
rect 562702 563378 588262 563614
rect 588498 563378 588670 563614
rect -4746 563366 588670 563378
rect -4746 563354 -4166 563366
rect 22294 563354 22874 563366
rect 58294 563354 58874 563366
rect 94294 563354 94874 563366
rect 130294 563354 130874 563366
rect 166294 563354 166874 563366
rect 202294 563354 202874 563366
rect 238294 563354 238874 563366
rect 274294 563354 274874 563366
rect 310294 563354 310874 563366
rect 346294 563354 346874 563366
rect 382294 563354 382874 563366
rect 418294 563354 418874 563366
rect 454294 563354 454874 563366
rect 490294 563354 490874 563366
rect 526294 563354 526874 563366
rect 562294 563354 562874 563366
rect 588090 563354 588670 563366
rect -2906 560466 -2326 560478
rect 18814 560466 19394 560478
rect 54814 560466 55394 560478
rect 90814 560466 91394 560478
rect 126814 560466 127394 560478
rect 162814 560466 163394 560478
rect 198814 560466 199394 560478
rect 234814 560466 235394 560478
rect 270814 560466 271394 560478
rect 306814 560466 307394 560478
rect 342814 560466 343394 560478
rect 378814 560466 379394 560478
rect 414814 560466 415394 560478
rect 450814 560466 451394 560478
rect 486814 560466 487394 560478
rect 522814 560466 523394 560478
rect 558814 560466 559394 560478
rect 586250 560466 586830 560478
rect -2906 560454 586830 560466
rect -2906 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586830 560454
rect -2906 560134 586830 560218
rect -2906 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586830 560134
rect -2906 559886 586830 559898
rect -2906 559874 -2326 559886
rect 18814 559874 19394 559886
rect 54814 559874 55394 559886
rect 90814 559874 91394 559886
rect 126814 559874 127394 559886
rect 162814 559874 163394 559886
rect 198814 559874 199394 559886
rect 234814 559874 235394 559886
rect 270814 559874 271394 559886
rect 306814 559874 307394 559886
rect 342814 559874 343394 559886
rect 378814 559874 379394 559886
rect 414814 559874 415394 559886
rect 450814 559874 451394 559886
rect 486814 559874 487394 559886
rect 522814 559874 523394 559886
rect 558814 559874 559394 559886
rect 586250 559874 586830 559886
rect -7506 552906 -6926 552918
rect 11254 552906 11834 552918
rect 47254 552906 47834 552918
rect 83254 552906 83834 552918
rect 119254 552906 119834 552918
rect 155254 552906 155834 552918
rect 191254 552906 191834 552918
rect 227254 552906 227834 552918
rect 263254 552906 263834 552918
rect 299254 552906 299834 552918
rect 335254 552906 335834 552918
rect 371254 552906 371834 552918
rect 407254 552906 407834 552918
rect 443254 552906 443834 552918
rect 479254 552906 479834 552918
rect 515254 552906 515834 552918
rect 551254 552906 551834 552918
rect 590850 552906 591430 552918
rect -8426 552894 592350 552906
rect -8426 552658 -7334 552894
rect -7098 552658 11426 552894
rect 11662 552658 47426 552894
rect 47662 552658 83426 552894
rect 83662 552658 119426 552894
rect 119662 552658 155426 552894
rect 155662 552658 191426 552894
rect 191662 552658 227426 552894
rect 227662 552658 263426 552894
rect 263662 552658 299426 552894
rect 299662 552658 335426 552894
rect 335662 552658 371426 552894
rect 371662 552658 407426 552894
rect 407662 552658 443426 552894
rect 443662 552658 479426 552894
rect 479662 552658 515426 552894
rect 515662 552658 551426 552894
rect 551662 552658 591022 552894
rect 591258 552658 592350 552894
rect -8426 552574 592350 552658
rect -8426 552338 -7334 552574
rect -7098 552338 11426 552574
rect 11662 552338 47426 552574
rect 47662 552338 83426 552574
rect 83662 552338 119426 552574
rect 119662 552338 155426 552574
rect 155662 552338 191426 552574
rect 191662 552338 227426 552574
rect 227662 552338 263426 552574
rect 263662 552338 299426 552574
rect 299662 552338 335426 552574
rect 335662 552338 371426 552574
rect 371662 552338 407426 552574
rect 407662 552338 443426 552574
rect 443662 552338 479426 552574
rect 479662 552338 515426 552574
rect 515662 552338 551426 552574
rect 551662 552338 591022 552574
rect 591258 552338 592350 552574
rect -8426 552326 592350 552338
rect -7506 552314 -6926 552326
rect 11254 552314 11834 552326
rect 47254 552314 47834 552326
rect 83254 552314 83834 552326
rect 119254 552314 119834 552326
rect 155254 552314 155834 552326
rect 191254 552314 191834 552326
rect 227254 552314 227834 552326
rect 263254 552314 263834 552326
rect 299254 552314 299834 552326
rect 335254 552314 335834 552326
rect 371254 552314 371834 552326
rect 407254 552314 407834 552326
rect 443254 552314 443834 552326
rect 479254 552314 479834 552326
rect 515254 552314 515834 552326
rect 551254 552314 551834 552326
rect 590850 552314 591430 552326
rect -5666 549426 -5086 549438
rect 7774 549426 8354 549438
rect 43774 549426 44354 549438
rect 79774 549426 80354 549438
rect 115774 549426 116354 549438
rect 151774 549426 152354 549438
rect 187774 549426 188354 549438
rect 223774 549426 224354 549438
rect 259774 549426 260354 549438
rect 295774 549426 296354 549438
rect 331774 549426 332354 549438
rect 367774 549426 368354 549438
rect 403774 549426 404354 549438
rect 439774 549426 440354 549438
rect 475774 549426 476354 549438
rect 511774 549426 512354 549438
rect 547774 549426 548354 549438
rect 589010 549426 589590 549438
rect -6586 549414 590510 549426
rect -6586 549178 -5494 549414
rect -5258 549178 7946 549414
rect 8182 549178 43946 549414
rect 44182 549178 79946 549414
rect 80182 549178 115946 549414
rect 116182 549178 151946 549414
rect 152182 549178 187946 549414
rect 188182 549178 223946 549414
rect 224182 549178 259946 549414
rect 260182 549178 295946 549414
rect 296182 549178 331946 549414
rect 332182 549178 367946 549414
rect 368182 549178 403946 549414
rect 404182 549178 439946 549414
rect 440182 549178 475946 549414
rect 476182 549178 511946 549414
rect 512182 549178 547946 549414
rect 548182 549178 589182 549414
rect 589418 549178 590510 549414
rect -6586 549094 590510 549178
rect -6586 548858 -5494 549094
rect -5258 548858 7946 549094
rect 8182 548858 43946 549094
rect 44182 548858 79946 549094
rect 80182 548858 115946 549094
rect 116182 548858 151946 549094
rect 152182 548858 187946 549094
rect 188182 548858 223946 549094
rect 224182 548858 259946 549094
rect 260182 548858 295946 549094
rect 296182 548858 331946 549094
rect 332182 548858 367946 549094
rect 368182 548858 403946 549094
rect 404182 548858 439946 549094
rect 440182 548858 475946 549094
rect 476182 548858 511946 549094
rect 512182 548858 547946 549094
rect 548182 548858 589182 549094
rect 589418 548858 590510 549094
rect -6586 548846 590510 548858
rect -5666 548834 -5086 548846
rect 7774 548834 8354 548846
rect 43774 548834 44354 548846
rect 79774 548834 80354 548846
rect 115774 548834 116354 548846
rect 151774 548834 152354 548846
rect 187774 548834 188354 548846
rect 223774 548834 224354 548846
rect 259774 548834 260354 548846
rect 295774 548834 296354 548846
rect 331774 548834 332354 548846
rect 367774 548834 368354 548846
rect 403774 548834 404354 548846
rect 439774 548834 440354 548846
rect 475774 548834 476354 548846
rect 511774 548834 512354 548846
rect 547774 548834 548354 548846
rect 589010 548834 589590 548846
rect -3826 545946 -3246 545958
rect 4294 545946 4874 545958
rect 40294 545946 40874 545958
rect 76294 545946 76874 545958
rect 112294 545946 112874 545958
rect 148294 545946 148874 545958
rect 184294 545946 184874 545958
rect 220294 545946 220874 545958
rect 256294 545946 256874 545958
rect 292294 545946 292874 545958
rect 328294 545946 328874 545958
rect 364294 545946 364874 545958
rect 400294 545946 400874 545958
rect 436294 545946 436874 545958
rect 472294 545946 472874 545958
rect 508294 545946 508874 545958
rect 544294 545946 544874 545958
rect 580294 545946 580874 545958
rect 587170 545946 587750 545958
rect -4746 545934 588670 545946
rect -4746 545698 -3654 545934
rect -3418 545698 4466 545934
rect 4702 545698 40466 545934
rect 40702 545698 76466 545934
rect 76702 545698 112466 545934
rect 112702 545698 148466 545934
rect 148702 545698 184466 545934
rect 184702 545698 220466 545934
rect 220702 545698 256466 545934
rect 256702 545698 292466 545934
rect 292702 545698 328466 545934
rect 328702 545698 364466 545934
rect 364702 545698 400466 545934
rect 400702 545698 436466 545934
rect 436702 545698 472466 545934
rect 472702 545698 508466 545934
rect 508702 545698 544466 545934
rect 544702 545698 580466 545934
rect 580702 545698 587342 545934
rect 587578 545698 588670 545934
rect -4746 545614 588670 545698
rect -4746 545378 -3654 545614
rect -3418 545378 4466 545614
rect 4702 545378 40466 545614
rect 40702 545378 76466 545614
rect 76702 545378 112466 545614
rect 112702 545378 148466 545614
rect 148702 545378 184466 545614
rect 184702 545378 220466 545614
rect 220702 545378 256466 545614
rect 256702 545378 292466 545614
rect 292702 545378 328466 545614
rect 328702 545378 364466 545614
rect 364702 545378 400466 545614
rect 400702 545378 436466 545614
rect 436702 545378 472466 545614
rect 472702 545378 508466 545614
rect 508702 545378 544466 545614
rect 544702 545378 580466 545614
rect 580702 545378 587342 545614
rect 587578 545378 588670 545614
rect -4746 545366 588670 545378
rect -3826 545354 -3246 545366
rect 4294 545354 4874 545366
rect 40294 545354 40874 545366
rect 76294 545354 76874 545366
rect 112294 545354 112874 545366
rect 148294 545354 148874 545366
rect 184294 545354 184874 545366
rect 220294 545354 220874 545366
rect 256294 545354 256874 545366
rect 292294 545354 292874 545366
rect 328294 545354 328874 545366
rect 364294 545354 364874 545366
rect 400294 545354 400874 545366
rect 436294 545354 436874 545366
rect 472294 545354 472874 545366
rect 508294 545354 508874 545366
rect 544294 545354 544874 545366
rect 580294 545354 580874 545366
rect 587170 545354 587750 545366
rect -1986 542466 -1406 542478
rect 814 542466 1394 542478
rect 36814 542466 37394 542478
rect 72814 542466 73394 542478
rect 108814 542466 109394 542478
rect 144814 542466 145394 542478
rect 180814 542466 181394 542478
rect 216814 542466 217394 542478
rect 252814 542466 253394 542478
rect 288814 542466 289394 542478
rect 324814 542466 325394 542478
rect 360814 542466 361394 542478
rect 396814 542466 397394 542478
rect 432814 542466 433394 542478
rect 468814 542466 469394 542478
rect 504814 542466 505394 542478
rect 540814 542466 541394 542478
rect 576814 542466 577394 542478
rect 585330 542466 585910 542478
rect -2906 542454 586830 542466
rect -2906 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586830 542454
rect -2906 542134 586830 542218
rect -2906 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586830 542134
rect -2906 541886 586830 541898
rect -1986 541874 -1406 541886
rect 814 541874 1394 541886
rect 36814 541874 37394 541886
rect 72814 541874 73394 541886
rect 108814 541874 109394 541886
rect 144814 541874 145394 541886
rect 180814 541874 181394 541886
rect 216814 541874 217394 541886
rect 252814 541874 253394 541886
rect 288814 541874 289394 541886
rect 324814 541874 325394 541886
rect 360814 541874 361394 541886
rect 396814 541874 397394 541886
rect 432814 541874 433394 541886
rect 468814 541874 469394 541886
rect 504814 541874 505394 541886
rect 540814 541874 541394 541886
rect 576814 541874 577394 541886
rect 585330 541874 585910 541886
rect -8426 534906 -7846 534918
rect 29254 534906 29834 534918
rect 65254 534906 65834 534918
rect 101254 534906 101834 534918
rect 137254 534906 137834 534918
rect 173254 534906 173834 534918
rect 209254 534906 209834 534918
rect 245254 534906 245834 534918
rect 281254 534906 281834 534918
rect 317254 534906 317834 534918
rect 353254 534906 353834 534918
rect 389254 534906 389834 534918
rect 425254 534906 425834 534918
rect 461254 534906 461834 534918
rect 497254 534906 497834 534918
rect 533254 534906 533834 534918
rect 569254 534906 569834 534918
rect 591770 534906 592350 534918
rect -8426 534894 592350 534906
rect -8426 534658 -8254 534894
rect -8018 534658 29426 534894
rect 29662 534658 65426 534894
rect 65662 534658 101426 534894
rect 101662 534658 137426 534894
rect 137662 534658 173426 534894
rect 173662 534658 209426 534894
rect 209662 534658 245426 534894
rect 245662 534658 281426 534894
rect 281662 534658 317426 534894
rect 317662 534658 353426 534894
rect 353662 534658 389426 534894
rect 389662 534658 425426 534894
rect 425662 534658 461426 534894
rect 461662 534658 497426 534894
rect 497662 534658 533426 534894
rect 533662 534658 569426 534894
rect 569662 534658 591942 534894
rect 592178 534658 592350 534894
rect -8426 534574 592350 534658
rect -8426 534338 -8254 534574
rect -8018 534338 29426 534574
rect 29662 534338 65426 534574
rect 65662 534338 101426 534574
rect 101662 534338 137426 534574
rect 137662 534338 173426 534574
rect 173662 534338 209426 534574
rect 209662 534338 245426 534574
rect 245662 534338 281426 534574
rect 281662 534338 317426 534574
rect 317662 534338 353426 534574
rect 353662 534338 389426 534574
rect 389662 534338 425426 534574
rect 425662 534338 461426 534574
rect 461662 534338 497426 534574
rect 497662 534338 533426 534574
rect 533662 534338 569426 534574
rect 569662 534338 591942 534574
rect 592178 534338 592350 534574
rect -8426 534326 592350 534338
rect -8426 534314 -7846 534326
rect 29254 534314 29834 534326
rect 65254 534314 65834 534326
rect 101254 534314 101834 534326
rect 137254 534314 137834 534326
rect 173254 534314 173834 534326
rect 209254 534314 209834 534326
rect 245254 534314 245834 534326
rect 281254 534314 281834 534326
rect 317254 534314 317834 534326
rect 353254 534314 353834 534326
rect 389254 534314 389834 534326
rect 425254 534314 425834 534326
rect 461254 534314 461834 534326
rect 497254 534314 497834 534326
rect 533254 534314 533834 534326
rect 569254 534314 569834 534326
rect 591770 534314 592350 534326
rect -6586 531426 -6006 531438
rect 25774 531426 26354 531438
rect 61774 531426 62354 531438
rect 97774 531426 98354 531438
rect 133774 531426 134354 531438
rect 169774 531426 170354 531438
rect 205774 531426 206354 531438
rect 241774 531426 242354 531438
rect 277774 531426 278354 531438
rect 313774 531426 314354 531438
rect 349774 531426 350354 531438
rect 385774 531426 386354 531438
rect 421774 531426 422354 531438
rect 457774 531426 458354 531438
rect 493774 531426 494354 531438
rect 529774 531426 530354 531438
rect 565774 531426 566354 531438
rect 589930 531426 590510 531438
rect -6586 531414 590510 531426
rect -6586 531178 -6414 531414
rect -6178 531178 25946 531414
rect 26182 531178 61946 531414
rect 62182 531178 97946 531414
rect 98182 531178 133946 531414
rect 134182 531178 169946 531414
rect 170182 531178 205946 531414
rect 206182 531178 241946 531414
rect 242182 531178 277946 531414
rect 278182 531178 313946 531414
rect 314182 531178 349946 531414
rect 350182 531178 385946 531414
rect 386182 531178 421946 531414
rect 422182 531178 457946 531414
rect 458182 531178 493946 531414
rect 494182 531178 529946 531414
rect 530182 531178 565946 531414
rect 566182 531178 590102 531414
rect 590338 531178 590510 531414
rect -6586 531094 590510 531178
rect -6586 530858 -6414 531094
rect -6178 530858 25946 531094
rect 26182 530858 61946 531094
rect 62182 530858 97946 531094
rect 98182 530858 133946 531094
rect 134182 530858 169946 531094
rect 170182 530858 205946 531094
rect 206182 530858 241946 531094
rect 242182 530858 277946 531094
rect 278182 530858 313946 531094
rect 314182 530858 349946 531094
rect 350182 530858 385946 531094
rect 386182 530858 421946 531094
rect 422182 530858 457946 531094
rect 458182 530858 493946 531094
rect 494182 530858 529946 531094
rect 530182 530858 565946 531094
rect 566182 530858 590102 531094
rect 590338 530858 590510 531094
rect -6586 530846 590510 530858
rect -6586 530834 -6006 530846
rect 25774 530834 26354 530846
rect 61774 530834 62354 530846
rect 97774 530834 98354 530846
rect 133774 530834 134354 530846
rect 169774 530834 170354 530846
rect 205774 530834 206354 530846
rect 241774 530834 242354 530846
rect 277774 530834 278354 530846
rect 313774 530834 314354 530846
rect 349774 530834 350354 530846
rect 385774 530834 386354 530846
rect 421774 530834 422354 530846
rect 457774 530834 458354 530846
rect 493774 530834 494354 530846
rect 529774 530834 530354 530846
rect 565774 530834 566354 530846
rect 589930 530834 590510 530846
rect -4746 527946 -4166 527958
rect 22294 527946 22874 527958
rect 58294 527946 58874 527958
rect 94294 527946 94874 527958
rect 130294 527946 130874 527958
rect 166294 527946 166874 527958
rect 202294 527946 202874 527958
rect 238294 527946 238874 527958
rect 274294 527946 274874 527958
rect 310294 527946 310874 527958
rect 346294 527946 346874 527958
rect 382294 527946 382874 527958
rect 418294 527946 418874 527958
rect 454294 527946 454874 527958
rect 490294 527946 490874 527958
rect 526294 527946 526874 527958
rect 562294 527946 562874 527958
rect 588090 527946 588670 527958
rect -4746 527934 588670 527946
rect -4746 527698 -4574 527934
rect -4338 527698 22466 527934
rect 22702 527698 58466 527934
rect 58702 527698 94466 527934
rect 94702 527698 130466 527934
rect 130702 527698 166466 527934
rect 166702 527698 202466 527934
rect 202702 527698 238466 527934
rect 238702 527698 274466 527934
rect 274702 527698 310466 527934
rect 310702 527698 346466 527934
rect 346702 527698 382466 527934
rect 382702 527698 418466 527934
rect 418702 527698 454466 527934
rect 454702 527698 490466 527934
rect 490702 527698 526466 527934
rect 526702 527698 562466 527934
rect 562702 527698 588262 527934
rect 588498 527698 588670 527934
rect -4746 527614 588670 527698
rect -4746 527378 -4574 527614
rect -4338 527378 22466 527614
rect 22702 527378 58466 527614
rect 58702 527378 94466 527614
rect 94702 527378 130466 527614
rect 130702 527378 166466 527614
rect 166702 527378 202466 527614
rect 202702 527378 238466 527614
rect 238702 527378 274466 527614
rect 274702 527378 310466 527614
rect 310702 527378 346466 527614
rect 346702 527378 382466 527614
rect 382702 527378 418466 527614
rect 418702 527378 454466 527614
rect 454702 527378 490466 527614
rect 490702 527378 526466 527614
rect 526702 527378 562466 527614
rect 562702 527378 588262 527614
rect 588498 527378 588670 527614
rect -4746 527366 588670 527378
rect -4746 527354 -4166 527366
rect 22294 527354 22874 527366
rect 58294 527354 58874 527366
rect 94294 527354 94874 527366
rect 130294 527354 130874 527366
rect 166294 527354 166874 527366
rect 202294 527354 202874 527366
rect 238294 527354 238874 527366
rect 274294 527354 274874 527366
rect 310294 527354 310874 527366
rect 346294 527354 346874 527366
rect 382294 527354 382874 527366
rect 418294 527354 418874 527366
rect 454294 527354 454874 527366
rect 490294 527354 490874 527366
rect 526294 527354 526874 527366
rect 562294 527354 562874 527366
rect 588090 527354 588670 527366
rect -2906 524466 -2326 524478
rect 18814 524466 19394 524478
rect 54814 524466 55394 524478
rect 90814 524466 91394 524478
rect 126814 524466 127394 524478
rect 162814 524466 163394 524478
rect 198814 524466 199394 524478
rect 234814 524466 235394 524478
rect 270814 524466 271394 524478
rect 306814 524466 307394 524478
rect 342814 524466 343394 524478
rect 378814 524466 379394 524478
rect 414814 524466 415394 524478
rect 450814 524466 451394 524478
rect 486814 524466 487394 524478
rect 522814 524466 523394 524478
rect 558814 524466 559394 524478
rect 586250 524466 586830 524478
rect -2906 524454 586830 524466
rect -2906 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586830 524454
rect -2906 524134 586830 524218
rect -2906 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586830 524134
rect -2906 523886 586830 523898
rect -2906 523874 -2326 523886
rect 18814 523874 19394 523886
rect 54814 523874 55394 523886
rect 90814 523874 91394 523886
rect 126814 523874 127394 523886
rect 162814 523874 163394 523886
rect 198814 523874 199394 523886
rect 234814 523874 235394 523886
rect 270814 523874 271394 523886
rect 306814 523874 307394 523886
rect 342814 523874 343394 523886
rect 378814 523874 379394 523886
rect 414814 523874 415394 523886
rect 450814 523874 451394 523886
rect 486814 523874 487394 523886
rect 522814 523874 523394 523886
rect 558814 523874 559394 523886
rect 586250 523874 586830 523886
rect -7506 516906 -6926 516918
rect 11254 516906 11834 516918
rect 47254 516906 47834 516918
rect 83254 516906 83834 516918
rect 119254 516906 119834 516918
rect 155254 516906 155834 516918
rect 191254 516906 191834 516918
rect 227254 516906 227834 516918
rect 263254 516906 263834 516918
rect 299254 516906 299834 516918
rect 335254 516906 335834 516918
rect 371254 516906 371834 516918
rect 407254 516906 407834 516918
rect 443254 516906 443834 516918
rect 479254 516906 479834 516918
rect 515254 516906 515834 516918
rect 551254 516906 551834 516918
rect 590850 516906 591430 516918
rect -8426 516894 592350 516906
rect -8426 516658 -7334 516894
rect -7098 516658 11426 516894
rect 11662 516658 47426 516894
rect 47662 516658 83426 516894
rect 83662 516658 119426 516894
rect 119662 516658 155426 516894
rect 155662 516658 191426 516894
rect 191662 516658 227426 516894
rect 227662 516658 263426 516894
rect 263662 516658 299426 516894
rect 299662 516658 335426 516894
rect 335662 516658 371426 516894
rect 371662 516658 407426 516894
rect 407662 516658 443426 516894
rect 443662 516658 479426 516894
rect 479662 516658 515426 516894
rect 515662 516658 551426 516894
rect 551662 516658 591022 516894
rect 591258 516658 592350 516894
rect -8426 516574 592350 516658
rect -8426 516338 -7334 516574
rect -7098 516338 11426 516574
rect 11662 516338 47426 516574
rect 47662 516338 83426 516574
rect 83662 516338 119426 516574
rect 119662 516338 155426 516574
rect 155662 516338 191426 516574
rect 191662 516338 227426 516574
rect 227662 516338 263426 516574
rect 263662 516338 299426 516574
rect 299662 516338 335426 516574
rect 335662 516338 371426 516574
rect 371662 516338 407426 516574
rect 407662 516338 443426 516574
rect 443662 516338 479426 516574
rect 479662 516338 515426 516574
rect 515662 516338 551426 516574
rect 551662 516338 591022 516574
rect 591258 516338 592350 516574
rect -8426 516326 592350 516338
rect -7506 516314 -6926 516326
rect 11254 516314 11834 516326
rect 47254 516314 47834 516326
rect 83254 516314 83834 516326
rect 119254 516314 119834 516326
rect 155254 516314 155834 516326
rect 191254 516314 191834 516326
rect 227254 516314 227834 516326
rect 263254 516314 263834 516326
rect 299254 516314 299834 516326
rect 335254 516314 335834 516326
rect 371254 516314 371834 516326
rect 407254 516314 407834 516326
rect 443254 516314 443834 516326
rect 479254 516314 479834 516326
rect 515254 516314 515834 516326
rect 551254 516314 551834 516326
rect 590850 516314 591430 516326
rect -5666 513426 -5086 513438
rect 7774 513426 8354 513438
rect 43774 513426 44354 513438
rect 79774 513426 80354 513438
rect 115774 513426 116354 513438
rect 151774 513426 152354 513438
rect 187774 513426 188354 513438
rect 223774 513426 224354 513438
rect 259774 513426 260354 513438
rect 295774 513426 296354 513438
rect 331774 513426 332354 513438
rect 367774 513426 368354 513438
rect 403774 513426 404354 513438
rect 439774 513426 440354 513438
rect 475774 513426 476354 513438
rect 511774 513426 512354 513438
rect 547774 513426 548354 513438
rect 589010 513426 589590 513438
rect -6586 513414 590510 513426
rect -6586 513178 -5494 513414
rect -5258 513178 7946 513414
rect 8182 513178 43946 513414
rect 44182 513178 79946 513414
rect 80182 513178 115946 513414
rect 116182 513178 151946 513414
rect 152182 513178 187946 513414
rect 188182 513178 223946 513414
rect 224182 513178 259946 513414
rect 260182 513178 295946 513414
rect 296182 513178 331946 513414
rect 332182 513178 367946 513414
rect 368182 513178 403946 513414
rect 404182 513178 439946 513414
rect 440182 513178 475946 513414
rect 476182 513178 511946 513414
rect 512182 513178 547946 513414
rect 548182 513178 589182 513414
rect 589418 513178 590510 513414
rect -6586 513094 590510 513178
rect -6586 512858 -5494 513094
rect -5258 512858 7946 513094
rect 8182 512858 43946 513094
rect 44182 512858 79946 513094
rect 80182 512858 115946 513094
rect 116182 512858 151946 513094
rect 152182 512858 187946 513094
rect 188182 512858 223946 513094
rect 224182 512858 259946 513094
rect 260182 512858 295946 513094
rect 296182 512858 331946 513094
rect 332182 512858 367946 513094
rect 368182 512858 403946 513094
rect 404182 512858 439946 513094
rect 440182 512858 475946 513094
rect 476182 512858 511946 513094
rect 512182 512858 547946 513094
rect 548182 512858 589182 513094
rect 589418 512858 590510 513094
rect -6586 512846 590510 512858
rect -5666 512834 -5086 512846
rect 7774 512834 8354 512846
rect 43774 512834 44354 512846
rect 79774 512834 80354 512846
rect 115774 512834 116354 512846
rect 151774 512834 152354 512846
rect 187774 512834 188354 512846
rect 223774 512834 224354 512846
rect 259774 512834 260354 512846
rect 295774 512834 296354 512846
rect 331774 512834 332354 512846
rect 367774 512834 368354 512846
rect 403774 512834 404354 512846
rect 439774 512834 440354 512846
rect 475774 512834 476354 512846
rect 511774 512834 512354 512846
rect 547774 512834 548354 512846
rect 589010 512834 589590 512846
rect -3826 509946 -3246 509958
rect 4294 509946 4874 509958
rect 40294 509946 40874 509958
rect 76294 509946 76874 509958
rect 112294 509946 112874 509958
rect 148294 509946 148874 509958
rect 184294 509946 184874 509958
rect 220294 509946 220874 509958
rect 256294 509946 256874 509958
rect 292294 509946 292874 509958
rect 328294 509946 328874 509958
rect 364294 509946 364874 509958
rect 400294 509946 400874 509958
rect 436294 509946 436874 509958
rect 472294 509946 472874 509958
rect 508294 509946 508874 509958
rect 544294 509946 544874 509958
rect 580294 509946 580874 509958
rect 587170 509946 587750 509958
rect -4746 509934 588670 509946
rect -4746 509698 -3654 509934
rect -3418 509698 4466 509934
rect 4702 509698 40466 509934
rect 40702 509698 76466 509934
rect 76702 509698 112466 509934
rect 112702 509698 148466 509934
rect 148702 509698 184466 509934
rect 184702 509698 220466 509934
rect 220702 509698 256466 509934
rect 256702 509698 292466 509934
rect 292702 509698 328466 509934
rect 328702 509698 364466 509934
rect 364702 509698 400466 509934
rect 400702 509698 436466 509934
rect 436702 509698 472466 509934
rect 472702 509698 508466 509934
rect 508702 509698 544466 509934
rect 544702 509698 580466 509934
rect 580702 509698 587342 509934
rect 587578 509698 588670 509934
rect -4746 509614 588670 509698
rect -4746 509378 -3654 509614
rect -3418 509378 4466 509614
rect 4702 509378 40466 509614
rect 40702 509378 76466 509614
rect 76702 509378 112466 509614
rect 112702 509378 148466 509614
rect 148702 509378 184466 509614
rect 184702 509378 220466 509614
rect 220702 509378 256466 509614
rect 256702 509378 292466 509614
rect 292702 509378 328466 509614
rect 328702 509378 364466 509614
rect 364702 509378 400466 509614
rect 400702 509378 436466 509614
rect 436702 509378 472466 509614
rect 472702 509378 508466 509614
rect 508702 509378 544466 509614
rect 544702 509378 580466 509614
rect 580702 509378 587342 509614
rect 587578 509378 588670 509614
rect -4746 509366 588670 509378
rect -3826 509354 -3246 509366
rect 4294 509354 4874 509366
rect 40294 509354 40874 509366
rect 76294 509354 76874 509366
rect 112294 509354 112874 509366
rect 148294 509354 148874 509366
rect 184294 509354 184874 509366
rect 220294 509354 220874 509366
rect 256294 509354 256874 509366
rect 292294 509354 292874 509366
rect 328294 509354 328874 509366
rect 364294 509354 364874 509366
rect 400294 509354 400874 509366
rect 436294 509354 436874 509366
rect 472294 509354 472874 509366
rect 508294 509354 508874 509366
rect 544294 509354 544874 509366
rect 580294 509354 580874 509366
rect 587170 509354 587750 509366
rect -1986 506466 -1406 506478
rect 814 506466 1394 506478
rect 36814 506466 37394 506478
rect 72814 506466 73394 506478
rect 108814 506466 109394 506478
rect 144814 506466 145394 506478
rect 180814 506466 181394 506478
rect 216814 506466 217394 506478
rect 252814 506466 253394 506478
rect 288814 506466 289394 506478
rect 324814 506466 325394 506478
rect 360814 506466 361394 506478
rect 396814 506466 397394 506478
rect 432814 506466 433394 506478
rect 468814 506466 469394 506478
rect 504814 506466 505394 506478
rect 540814 506466 541394 506478
rect 576814 506466 577394 506478
rect 585330 506466 585910 506478
rect -2906 506454 586830 506466
rect -2906 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586830 506454
rect -2906 506134 586830 506218
rect -2906 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586830 506134
rect -2906 505886 586830 505898
rect -1986 505874 -1406 505886
rect 814 505874 1394 505886
rect 36814 505874 37394 505886
rect 72814 505874 73394 505886
rect 108814 505874 109394 505886
rect 144814 505874 145394 505886
rect 180814 505874 181394 505886
rect 216814 505874 217394 505886
rect 252814 505874 253394 505886
rect 288814 505874 289394 505886
rect 324814 505874 325394 505886
rect 360814 505874 361394 505886
rect 396814 505874 397394 505886
rect 432814 505874 433394 505886
rect 468814 505874 469394 505886
rect 504814 505874 505394 505886
rect 540814 505874 541394 505886
rect 576814 505874 577394 505886
rect 585330 505874 585910 505886
rect -8426 498906 -7846 498918
rect 29254 498906 29834 498918
rect 65254 498906 65834 498918
rect 101254 498906 101834 498918
rect 137254 498906 137834 498918
rect 173254 498906 173834 498918
rect 209254 498906 209834 498918
rect 245254 498906 245834 498918
rect 281254 498906 281834 498918
rect 317254 498906 317834 498918
rect 353254 498906 353834 498918
rect 389254 498906 389834 498918
rect 425254 498906 425834 498918
rect 461254 498906 461834 498918
rect 497254 498906 497834 498918
rect 533254 498906 533834 498918
rect 569254 498906 569834 498918
rect 591770 498906 592350 498918
rect -8426 498894 592350 498906
rect -8426 498658 -8254 498894
rect -8018 498658 29426 498894
rect 29662 498658 65426 498894
rect 65662 498658 101426 498894
rect 101662 498658 137426 498894
rect 137662 498658 173426 498894
rect 173662 498658 209426 498894
rect 209662 498658 245426 498894
rect 245662 498658 281426 498894
rect 281662 498658 317426 498894
rect 317662 498658 353426 498894
rect 353662 498658 389426 498894
rect 389662 498658 425426 498894
rect 425662 498658 461426 498894
rect 461662 498658 497426 498894
rect 497662 498658 533426 498894
rect 533662 498658 569426 498894
rect 569662 498658 591942 498894
rect 592178 498658 592350 498894
rect -8426 498574 592350 498658
rect -8426 498338 -8254 498574
rect -8018 498338 29426 498574
rect 29662 498338 65426 498574
rect 65662 498338 101426 498574
rect 101662 498338 137426 498574
rect 137662 498338 173426 498574
rect 173662 498338 209426 498574
rect 209662 498338 245426 498574
rect 245662 498338 281426 498574
rect 281662 498338 317426 498574
rect 317662 498338 353426 498574
rect 353662 498338 389426 498574
rect 389662 498338 425426 498574
rect 425662 498338 461426 498574
rect 461662 498338 497426 498574
rect 497662 498338 533426 498574
rect 533662 498338 569426 498574
rect 569662 498338 591942 498574
rect 592178 498338 592350 498574
rect -8426 498326 592350 498338
rect -8426 498314 -7846 498326
rect 29254 498314 29834 498326
rect 65254 498314 65834 498326
rect 101254 498314 101834 498326
rect 137254 498314 137834 498326
rect 173254 498314 173834 498326
rect 209254 498314 209834 498326
rect 245254 498314 245834 498326
rect 281254 498314 281834 498326
rect 317254 498314 317834 498326
rect 353254 498314 353834 498326
rect 389254 498314 389834 498326
rect 425254 498314 425834 498326
rect 461254 498314 461834 498326
rect 497254 498314 497834 498326
rect 533254 498314 533834 498326
rect 569254 498314 569834 498326
rect 591770 498314 592350 498326
rect -6586 495426 -6006 495438
rect 25774 495426 26354 495438
rect 61774 495426 62354 495438
rect 97774 495426 98354 495438
rect 133774 495426 134354 495438
rect 169774 495426 170354 495438
rect 205774 495426 206354 495438
rect 241774 495426 242354 495438
rect 277774 495426 278354 495438
rect 313774 495426 314354 495438
rect 349774 495426 350354 495438
rect 385774 495426 386354 495438
rect 421774 495426 422354 495438
rect 457774 495426 458354 495438
rect 493774 495426 494354 495438
rect 529774 495426 530354 495438
rect 565774 495426 566354 495438
rect 589930 495426 590510 495438
rect -6586 495414 590510 495426
rect -6586 495178 -6414 495414
rect -6178 495178 25946 495414
rect 26182 495178 61946 495414
rect 62182 495178 97946 495414
rect 98182 495178 133946 495414
rect 134182 495178 169946 495414
rect 170182 495178 205946 495414
rect 206182 495178 241946 495414
rect 242182 495178 277946 495414
rect 278182 495178 313946 495414
rect 314182 495178 349946 495414
rect 350182 495178 385946 495414
rect 386182 495178 421946 495414
rect 422182 495178 457946 495414
rect 458182 495178 493946 495414
rect 494182 495178 529946 495414
rect 530182 495178 565946 495414
rect 566182 495178 590102 495414
rect 590338 495178 590510 495414
rect -6586 495094 590510 495178
rect -6586 494858 -6414 495094
rect -6178 494858 25946 495094
rect 26182 494858 61946 495094
rect 62182 494858 97946 495094
rect 98182 494858 133946 495094
rect 134182 494858 169946 495094
rect 170182 494858 205946 495094
rect 206182 494858 241946 495094
rect 242182 494858 277946 495094
rect 278182 494858 313946 495094
rect 314182 494858 349946 495094
rect 350182 494858 385946 495094
rect 386182 494858 421946 495094
rect 422182 494858 457946 495094
rect 458182 494858 493946 495094
rect 494182 494858 529946 495094
rect 530182 494858 565946 495094
rect 566182 494858 590102 495094
rect 590338 494858 590510 495094
rect -6586 494846 590510 494858
rect -6586 494834 -6006 494846
rect 25774 494834 26354 494846
rect 61774 494834 62354 494846
rect 97774 494834 98354 494846
rect 133774 494834 134354 494846
rect 169774 494834 170354 494846
rect 205774 494834 206354 494846
rect 241774 494834 242354 494846
rect 277774 494834 278354 494846
rect 313774 494834 314354 494846
rect 349774 494834 350354 494846
rect 385774 494834 386354 494846
rect 421774 494834 422354 494846
rect 457774 494834 458354 494846
rect 493774 494834 494354 494846
rect 529774 494834 530354 494846
rect 565774 494834 566354 494846
rect 589930 494834 590510 494846
rect -4746 491946 -4166 491958
rect 22294 491946 22874 491958
rect 58294 491946 58874 491958
rect 94294 491946 94874 491958
rect 130294 491946 130874 491958
rect 166294 491946 166874 491958
rect 202294 491946 202874 491958
rect 238294 491946 238874 491958
rect 274294 491946 274874 491958
rect 310294 491946 310874 491958
rect 346294 491946 346874 491958
rect 382294 491946 382874 491958
rect 418294 491946 418874 491958
rect 454294 491946 454874 491958
rect 490294 491946 490874 491958
rect 526294 491946 526874 491958
rect 562294 491946 562874 491958
rect 588090 491946 588670 491958
rect -4746 491934 588670 491946
rect -4746 491698 -4574 491934
rect -4338 491698 22466 491934
rect 22702 491698 58466 491934
rect 58702 491698 94466 491934
rect 94702 491698 130466 491934
rect 130702 491698 166466 491934
rect 166702 491698 202466 491934
rect 202702 491698 238466 491934
rect 238702 491698 274466 491934
rect 274702 491698 310466 491934
rect 310702 491698 346466 491934
rect 346702 491698 382466 491934
rect 382702 491698 418466 491934
rect 418702 491698 454466 491934
rect 454702 491698 490466 491934
rect 490702 491698 526466 491934
rect 526702 491698 562466 491934
rect 562702 491698 588262 491934
rect 588498 491698 588670 491934
rect -4746 491614 588670 491698
rect -4746 491378 -4574 491614
rect -4338 491378 22466 491614
rect 22702 491378 58466 491614
rect 58702 491378 94466 491614
rect 94702 491378 130466 491614
rect 130702 491378 166466 491614
rect 166702 491378 202466 491614
rect 202702 491378 238466 491614
rect 238702 491378 274466 491614
rect 274702 491378 310466 491614
rect 310702 491378 346466 491614
rect 346702 491378 382466 491614
rect 382702 491378 418466 491614
rect 418702 491378 454466 491614
rect 454702 491378 490466 491614
rect 490702 491378 526466 491614
rect 526702 491378 562466 491614
rect 562702 491378 588262 491614
rect 588498 491378 588670 491614
rect -4746 491366 588670 491378
rect -4746 491354 -4166 491366
rect 22294 491354 22874 491366
rect 58294 491354 58874 491366
rect 94294 491354 94874 491366
rect 130294 491354 130874 491366
rect 166294 491354 166874 491366
rect 202294 491354 202874 491366
rect 238294 491354 238874 491366
rect 274294 491354 274874 491366
rect 310294 491354 310874 491366
rect 346294 491354 346874 491366
rect 382294 491354 382874 491366
rect 418294 491354 418874 491366
rect 454294 491354 454874 491366
rect 490294 491354 490874 491366
rect 526294 491354 526874 491366
rect 562294 491354 562874 491366
rect 588090 491354 588670 491366
rect -2906 488466 -2326 488478
rect 18814 488466 19394 488478
rect 54814 488466 55394 488478
rect 90814 488466 91394 488478
rect 126814 488466 127394 488478
rect 162814 488466 163394 488478
rect 198814 488466 199394 488478
rect 234814 488466 235394 488478
rect 270814 488466 271394 488478
rect 306814 488466 307394 488478
rect 342814 488466 343394 488478
rect 378814 488466 379394 488478
rect 414814 488466 415394 488478
rect 450814 488466 451394 488478
rect 486814 488466 487394 488478
rect 522814 488466 523394 488478
rect 558814 488466 559394 488478
rect 586250 488466 586830 488478
rect -2906 488454 586830 488466
rect -2906 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586830 488454
rect -2906 488134 586830 488218
rect -2906 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586830 488134
rect -2906 487886 586830 487898
rect -2906 487874 -2326 487886
rect 18814 487874 19394 487886
rect 54814 487874 55394 487886
rect 90814 487874 91394 487886
rect 126814 487874 127394 487886
rect 162814 487874 163394 487886
rect 198814 487874 199394 487886
rect 234814 487874 235394 487886
rect 270814 487874 271394 487886
rect 306814 487874 307394 487886
rect 342814 487874 343394 487886
rect 378814 487874 379394 487886
rect 414814 487874 415394 487886
rect 450814 487874 451394 487886
rect 486814 487874 487394 487886
rect 522814 487874 523394 487886
rect 558814 487874 559394 487886
rect 586250 487874 586830 487886
rect -7506 480906 -6926 480918
rect 11254 480906 11834 480918
rect 47254 480906 47834 480918
rect 83254 480906 83834 480918
rect 119254 480906 119834 480918
rect 155254 480906 155834 480918
rect 191254 480906 191834 480918
rect 227254 480906 227834 480918
rect 263254 480906 263834 480918
rect 299254 480906 299834 480918
rect 335254 480906 335834 480918
rect 371254 480906 371834 480918
rect 407254 480906 407834 480918
rect 443254 480906 443834 480918
rect 479254 480906 479834 480918
rect 515254 480906 515834 480918
rect 551254 480906 551834 480918
rect 590850 480906 591430 480918
rect -8426 480894 592350 480906
rect -8426 480658 -7334 480894
rect -7098 480658 11426 480894
rect 11662 480658 47426 480894
rect 47662 480658 83426 480894
rect 83662 480658 119426 480894
rect 119662 480658 155426 480894
rect 155662 480658 191426 480894
rect 191662 480658 227426 480894
rect 227662 480658 263426 480894
rect 263662 480658 299426 480894
rect 299662 480658 335426 480894
rect 335662 480658 371426 480894
rect 371662 480658 407426 480894
rect 407662 480658 443426 480894
rect 443662 480658 479426 480894
rect 479662 480658 515426 480894
rect 515662 480658 551426 480894
rect 551662 480658 591022 480894
rect 591258 480658 592350 480894
rect -8426 480574 592350 480658
rect -8426 480338 -7334 480574
rect -7098 480338 11426 480574
rect 11662 480338 47426 480574
rect 47662 480338 83426 480574
rect 83662 480338 119426 480574
rect 119662 480338 155426 480574
rect 155662 480338 191426 480574
rect 191662 480338 227426 480574
rect 227662 480338 263426 480574
rect 263662 480338 299426 480574
rect 299662 480338 335426 480574
rect 335662 480338 371426 480574
rect 371662 480338 407426 480574
rect 407662 480338 443426 480574
rect 443662 480338 479426 480574
rect 479662 480338 515426 480574
rect 515662 480338 551426 480574
rect 551662 480338 591022 480574
rect 591258 480338 592350 480574
rect -8426 480326 592350 480338
rect -7506 480314 -6926 480326
rect 11254 480314 11834 480326
rect 47254 480314 47834 480326
rect 83254 480314 83834 480326
rect 119254 480314 119834 480326
rect 155254 480314 155834 480326
rect 191254 480314 191834 480326
rect 227254 480314 227834 480326
rect 263254 480314 263834 480326
rect 299254 480314 299834 480326
rect 335254 480314 335834 480326
rect 371254 480314 371834 480326
rect 407254 480314 407834 480326
rect 443254 480314 443834 480326
rect 479254 480314 479834 480326
rect 515254 480314 515834 480326
rect 551254 480314 551834 480326
rect 590850 480314 591430 480326
rect -5666 477426 -5086 477438
rect 7774 477426 8354 477438
rect 43774 477426 44354 477438
rect 79774 477426 80354 477438
rect 115774 477426 116354 477438
rect 151774 477426 152354 477438
rect 187774 477426 188354 477438
rect 223774 477426 224354 477438
rect 259774 477426 260354 477438
rect 295774 477426 296354 477438
rect 331774 477426 332354 477438
rect 367774 477426 368354 477438
rect 403774 477426 404354 477438
rect 439774 477426 440354 477438
rect 475774 477426 476354 477438
rect 511774 477426 512354 477438
rect 547774 477426 548354 477438
rect 589010 477426 589590 477438
rect -6586 477414 590510 477426
rect -6586 477178 -5494 477414
rect -5258 477178 7946 477414
rect 8182 477178 43946 477414
rect 44182 477178 79946 477414
rect 80182 477178 115946 477414
rect 116182 477178 151946 477414
rect 152182 477178 187946 477414
rect 188182 477178 223946 477414
rect 224182 477178 259946 477414
rect 260182 477178 295946 477414
rect 296182 477178 331946 477414
rect 332182 477178 367946 477414
rect 368182 477178 403946 477414
rect 404182 477178 439946 477414
rect 440182 477178 475946 477414
rect 476182 477178 511946 477414
rect 512182 477178 547946 477414
rect 548182 477178 589182 477414
rect 589418 477178 590510 477414
rect -6586 477094 590510 477178
rect -6586 476858 -5494 477094
rect -5258 476858 7946 477094
rect 8182 476858 43946 477094
rect 44182 476858 79946 477094
rect 80182 476858 115946 477094
rect 116182 476858 151946 477094
rect 152182 476858 187946 477094
rect 188182 476858 223946 477094
rect 224182 476858 259946 477094
rect 260182 476858 295946 477094
rect 296182 476858 331946 477094
rect 332182 476858 367946 477094
rect 368182 476858 403946 477094
rect 404182 476858 439946 477094
rect 440182 476858 475946 477094
rect 476182 476858 511946 477094
rect 512182 476858 547946 477094
rect 548182 476858 589182 477094
rect 589418 476858 590510 477094
rect -6586 476846 590510 476858
rect -5666 476834 -5086 476846
rect 7774 476834 8354 476846
rect 43774 476834 44354 476846
rect 79774 476834 80354 476846
rect 115774 476834 116354 476846
rect 151774 476834 152354 476846
rect 187774 476834 188354 476846
rect 223774 476834 224354 476846
rect 259774 476834 260354 476846
rect 295774 476834 296354 476846
rect 331774 476834 332354 476846
rect 367774 476834 368354 476846
rect 403774 476834 404354 476846
rect 439774 476834 440354 476846
rect 475774 476834 476354 476846
rect 511774 476834 512354 476846
rect 547774 476834 548354 476846
rect 589010 476834 589590 476846
rect -3826 473946 -3246 473958
rect 4294 473946 4874 473958
rect 40294 473946 40874 473958
rect 76294 473946 76874 473958
rect 112294 473946 112874 473958
rect 148294 473946 148874 473958
rect 184294 473946 184874 473958
rect 220294 473946 220874 473958
rect 256294 473946 256874 473958
rect 292294 473946 292874 473958
rect 328294 473946 328874 473958
rect 364294 473946 364874 473958
rect 400294 473946 400874 473958
rect 436294 473946 436874 473958
rect 472294 473946 472874 473958
rect 508294 473946 508874 473958
rect 544294 473946 544874 473958
rect 580294 473946 580874 473958
rect 587170 473946 587750 473958
rect -4746 473934 588670 473946
rect -4746 473698 -3654 473934
rect -3418 473698 4466 473934
rect 4702 473698 40466 473934
rect 40702 473698 76466 473934
rect 76702 473698 112466 473934
rect 112702 473698 148466 473934
rect 148702 473698 184466 473934
rect 184702 473698 220466 473934
rect 220702 473698 256466 473934
rect 256702 473698 292466 473934
rect 292702 473698 328466 473934
rect 328702 473698 364466 473934
rect 364702 473698 400466 473934
rect 400702 473698 436466 473934
rect 436702 473698 472466 473934
rect 472702 473698 508466 473934
rect 508702 473698 544466 473934
rect 544702 473698 580466 473934
rect 580702 473698 587342 473934
rect 587578 473698 588670 473934
rect -4746 473614 588670 473698
rect -4746 473378 -3654 473614
rect -3418 473378 4466 473614
rect 4702 473378 40466 473614
rect 40702 473378 76466 473614
rect 76702 473378 112466 473614
rect 112702 473378 148466 473614
rect 148702 473378 184466 473614
rect 184702 473378 220466 473614
rect 220702 473378 256466 473614
rect 256702 473378 292466 473614
rect 292702 473378 328466 473614
rect 328702 473378 364466 473614
rect 364702 473378 400466 473614
rect 400702 473378 436466 473614
rect 436702 473378 472466 473614
rect 472702 473378 508466 473614
rect 508702 473378 544466 473614
rect 544702 473378 580466 473614
rect 580702 473378 587342 473614
rect 587578 473378 588670 473614
rect -4746 473366 588670 473378
rect -3826 473354 -3246 473366
rect 4294 473354 4874 473366
rect 40294 473354 40874 473366
rect 76294 473354 76874 473366
rect 112294 473354 112874 473366
rect 148294 473354 148874 473366
rect 184294 473354 184874 473366
rect 220294 473354 220874 473366
rect 256294 473354 256874 473366
rect 292294 473354 292874 473366
rect 328294 473354 328874 473366
rect 364294 473354 364874 473366
rect 400294 473354 400874 473366
rect 436294 473354 436874 473366
rect 472294 473354 472874 473366
rect 508294 473354 508874 473366
rect 544294 473354 544874 473366
rect 580294 473354 580874 473366
rect 587170 473354 587750 473366
rect -1986 470466 -1406 470478
rect 814 470466 1394 470478
rect 36814 470466 37394 470478
rect 72814 470466 73394 470478
rect 108814 470466 109394 470478
rect 144814 470466 145394 470478
rect 180814 470466 181394 470478
rect 216814 470466 217394 470478
rect 252814 470466 253394 470478
rect 288814 470466 289394 470478
rect 324814 470466 325394 470478
rect 360814 470466 361394 470478
rect 396814 470466 397394 470478
rect 432814 470466 433394 470478
rect 468814 470466 469394 470478
rect 504814 470466 505394 470478
rect 540814 470466 541394 470478
rect 576814 470466 577394 470478
rect 585330 470466 585910 470478
rect -2906 470454 586830 470466
rect -2906 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586830 470454
rect -2906 470134 586830 470218
rect -2906 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586830 470134
rect -2906 469886 586830 469898
rect -1986 469874 -1406 469886
rect 814 469874 1394 469886
rect 36814 469874 37394 469886
rect 72814 469874 73394 469886
rect 108814 469874 109394 469886
rect 144814 469874 145394 469886
rect 180814 469874 181394 469886
rect 216814 469874 217394 469886
rect 252814 469874 253394 469886
rect 288814 469874 289394 469886
rect 324814 469874 325394 469886
rect 360814 469874 361394 469886
rect 396814 469874 397394 469886
rect 432814 469874 433394 469886
rect 468814 469874 469394 469886
rect 504814 469874 505394 469886
rect 540814 469874 541394 469886
rect 576814 469874 577394 469886
rect 585330 469874 585910 469886
rect -8426 462906 -7846 462918
rect 29254 462906 29834 462918
rect 65254 462906 65834 462918
rect 101254 462906 101834 462918
rect 137254 462906 137834 462918
rect 173254 462906 173834 462918
rect 209254 462906 209834 462918
rect 245254 462906 245834 462918
rect 281254 462906 281834 462918
rect 317254 462906 317834 462918
rect 353254 462906 353834 462918
rect 389254 462906 389834 462918
rect 425254 462906 425834 462918
rect 461254 462906 461834 462918
rect 497254 462906 497834 462918
rect 533254 462906 533834 462918
rect 569254 462906 569834 462918
rect 591770 462906 592350 462918
rect -8426 462894 592350 462906
rect -8426 462658 -8254 462894
rect -8018 462658 29426 462894
rect 29662 462658 65426 462894
rect 65662 462658 101426 462894
rect 101662 462658 137426 462894
rect 137662 462658 173426 462894
rect 173662 462658 209426 462894
rect 209662 462658 245426 462894
rect 245662 462658 281426 462894
rect 281662 462658 317426 462894
rect 317662 462658 353426 462894
rect 353662 462658 389426 462894
rect 389662 462658 425426 462894
rect 425662 462658 461426 462894
rect 461662 462658 497426 462894
rect 497662 462658 533426 462894
rect 533662 462658 569426 462894
rect 569662 462658 591942 462894
rect 592178 462658 592350 462894
rect -8426 462574 592350 462658
rect -8426 462338 -8254 462574
rect -8018 462338 29426 462574
rect 29662 462338 65426 462574
rect 65662 462338 101426 462574
rect 101662 462338 137426 462574
rect 137662 462338 173426 462574
rect 173662 462338 209426 462574
rect 209662 462338 245426 462574
rect 245662 462338 281426 462574
rect 281662 462338 317426 462574
rect 317662 462338 353426 462574
rect 353662 462338 389426 462574
rect 389662 462338 425426 462574
rect 425662 462338 461426 462574
rect 461662 462338 497426 462574
rect 497662 462338 533426 462574
rect 533662 462338 569426 462574
rect 569662 462338 591942 462574
rect 592178 462338 592350 462574
rect -8426 462326 592350 462338
rect -8426 462314 -7846 462326
rect 29254 462314 29834 462326
rect 65254 462314 65834 462326
rect 101254 462314 101834 462326
rect 137254 462314 137834 462326
rect 173254 462314 173834 462326
rect 209254 462314 209834 462326
rect 245254 462314 245834 462326
rect 281254 462314 281834 462326
rect 317254 462314 317834 462326
rect 353254 462314 353834 462326
rect 389254 462314 389834 462326
rect 425254 462314 425834 462326
rect 461254 462314 461834 462326
rect 497254 462314 497834 462326
rect 533254 462314 533834 462326
rect 569254 462314 569834 462326
rect 591770 462314 592350 462326
rect -6586 459426 -6006 459438
rect 25774 459426 26354 459438
rect 61774 459426 62354 459438
rect 97774 459426 98354 459438
rect 133774 459426 134354 459438
rect 169774 459426 170354 459438
rect 205774 459426 206354 459438
rect 241774 459426 242354 459438
rect 277774 459426 278354 459438
rect 313774 459426 314354 459438
rect 349774 459426 350354 459438
rect 385774 459426 386354 459438
rect 421774 459426 422354 459438
rect 457774 459426 458354 459438
rect 493774 459426 494354 459438
rect 529774 459426 530354 459438
rect 565774 459426 566354 459438
rect 589930 459426 590510 459438
rect -6586 459414 590510 459426
rect -6586 459178 -6414 459414
rect -6178 459178 25946 459414
rect 26182 459178 61946 459414
rect 62182 459178 97946 459414
rect 98182 459178 133946 459414
rect 134182 459178 169946 459414
rect 170182 459178 205946 459414
rect 206182 459178 241946 459414
rect 242182 459178 277946 459414
rect 278182 459178 313946 459414
rect 314182 459178 349946 459414
rect 350182 459178 385946 459414
rect 386182 459178 421946 459414
rect 422182 459178 457946 459414
rect 458182 459178 493946 459414
rect 494182 459178 529946 459414
rect 530182 459178 565946 459414
rect 566182 459178 590102 459414
rect 590338 459178 590510 459414
rect -6586 459094 590510 459178
rect -6586 458858 -6414 459094
rect -6178 458858 25946 459094
rect 26182 458858 61946 459094
rect 62182 458858 97946 459094
rect 98182 458858 133946 459094
rect 134182 458858 169946 459094
rect 170182 458858 205946 459094
rect 206182 458858 241946 459094
rect 242182 458858 277946 459094
rect 278182 458858 313946 459094
rect 314182 458858 349946 459094
rect 350182 458858 385946 459094
rect 386182 458858 421946 459094
rect 422182 458858 457946 459094
rect 458182 458858 493946 459094
rect 494182 458858 529946 459094
rect 530182 458858 565946 459094
rect 566182 458858 590102 459094
rect 590338 458858 590510 459094
rect -6586 458846 590510 458858
rect -6586 458834 -6006 458846
rect 25774 458834 26354 458846
rect 61774 458834 62354 458846
rect 97774 458834 98354 458846
rect 133774 458834 134354 458846
rect 169774 458834 170354 458846
rect 205774 458834 206354 458846
rect 241774 458834 242354 458846
rect 277774 458834 278354 458846
rect 313774 458834 314354 458846
rect 349774 458834 350354 458846
rect 385774 458834 386354 458846
rect 421774 458834 422354 458846
rect 457774 458834 458354 458846
rect 493774 458834 494354 458846
rect 529774 458834 530354 458846
rect 565774 458834 566354 458846
rect 589930 458834 590510 458846
rect -4746 455946 -4166 455958
rect 22294 455946 22874 455958
rect 58294 455946 58874 455958
rect 94294 455946 94874 455958
rect 130294 455946 130874 455958
rect 166294 455946 166874 455958
rect 202294 455946 202874 455958
rect 238294 455946 238874 455958
rect 274294 455946 274874 455958
rect 310294 455946 310874 455958
rect 346294 455946 346874 455958
rect 382294 455946 382874 455958
rect 418294 455946 418874 455958
rect 454294 455946 454874 455958
rect 490294 455946 490874 455958
rect 526294 455946 526874 455958
rect 562294 455946 562874 455958
rect 588090 455946 588670 455958
rect -4746 455934 588670 455946
rect -4746 455698 -4574 455934
rect -4338 455698 22466 455934
rect 22702 455698 58466 455934
rect 58702 455698 94466 455934
rect 94702 455698 130466 455934
rect 130702 455698 166466 455934
rect 166702 455698 202466 455934
rect 202702 455698 238466 455934
rect 238702 455698 274466 455934
rect 274702 455698 310466 455934
rect 310702 455698 346466 455934
rect 346702 455698 382466 455934
rect 382702 455698 418466 455934
rect 418702 455698 454466 455934
rect 454702 455698 490466 455934
rect 490702 455698 526466 455934
rect 526702 455698 562466 455934
rect 562702 455698 588262 455934
rect 588498 455698 588670 455934
rect -4746 455614 588670 455698
rect -4746 455378 -4574 455614
rect -4338 455378 22466 455614
rect 22702 455378 58466 455614
rect 58702 455378 94466 455614
rect 94702 455378 130466 455614
rect 130702 455378 166466 455614
rect 166702 455378 202466 455614
rect 202702 455378 238466 455614
rect 238702 455378 274466 455614
rect 274702 455378 310466 455614
rect 310702 455378 346466 455614
rect 346702 455378 382466 455614
rect 382702 455378 418466 455614
rect 418702 455378 454466 455614
rect 454702 455378 490466 455614
rect 490702 455378 526466 455614
rect 526702 455378 562466 455614
rect 562702 455378 588262 455614
rect 588498 455378 588670 455614
rect -4746 455366 588670 455378
rect -4746 455354 -4166 455366
rect 22294 455354 22874 455366
rect 58294 455354 58874 455366
rect 94294 455354 94874 455366
rect 130294 455354 130874 455366
rect 166294 455354 166874 455366
rect 202294 455354 202874 455366
rect 238294 455354 238874 455366
rect 274294 455354 274874 455366
rect 310294 455354 310874 455366
rect 346294 455354 346874 455366
rect 382294 455354 382874 455366
rect 418294 455354 418874 455366
rect 454294 455354 454874 455366
rect 490294 455354 490874 455366
rect 526294 455354 526874 455366
rect 562294 455354 562874 455366
rect 588090 455354 588670 455366
rect -2906 452466 -2326 452478
rect 18814 452466 19394 452478
rect 54814 452466 55394 452478
rect 90814 452466 91394 452478
rect 126814 452466 127394 452478
rect 162814 452466 163394 452478
rect 198814 452466 199394 452478
rect 234814 452466 235394 452478
rect 270814 452466 271394 452478
rect 306814 452466 307394 452478
rect 342814 452466 343394 452478
rect 378814 452466 379394 452478
rect 414814 452466 415394 452478
rect 450814 452466 451394 452478
rect 486814 452466 487394 452478
rect 522814 452466 523394 452478
rect 558814 452466 559394 452478
rect 586250 452466 586830 452478
rect -2906 452454 586830 452466
rect -2906 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586830 452454
rect -2906 452134 586830 452218
rect -2906 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586830 452134
rect -2906 451886 586830 451898
rect -2906 451874 -2326 451886
rect 18814 451874 19394 451886
rect 54814 451874 55394 451886
rect 90814 451874 91394 451886
rect 126814 451874 127394 451886
rect 162814 451874 163394 451886
rect 198814 451874 199394 451886
rect 234814 451874 235394 451886
rect 270814 451874 271394 451886
rect 306814 451874 307394 451886
rect 342814 451874 343394 451886
rect 378814 451874 379394 451886
rect 414814 451874 415394 451886
rect 450814 451874 451394 451886
rect 486814 451874 487394 451886
rect 522814 451874 523394 451886
rect 558814 451874 559394 451886
rect 586250 451874 586830 451886
rect -7506 444906 -6926 444918
rect 11254 444906 11834 444918
rect 47254 444906 47834 444918
rect 83254 444906 83834 444918
rect 119254 444906 119834 444918
rect 155254 444906 155834 444918
rect 191254 444906 191834 444918
rect 227254 444906 227834 444918
rect 263254 444906 263834 444918
rect 299254 444906 299834 444918
rect 335254 444906 335834 444918
rect 371254 444906 371834 444918
rect 407254 444906 407834 444918
rect 443254 444906 443834 444918
rect 479254 444906 479834 444918
rect 515254 444906 515834 444918
rect 551254 444906 551834 444918
rect 590850 444906 591430 444918
rect -8426 444894 592350 444906
rect -8426 444658 -7334 444894
rect -7098 444658 11426 444894
rect 11662 444658 47426 444894
rect 47662 444658 83426 444894
rect 83662 444658 119426 444894
rect 119662 444658 155426 444894
rect 155662 444658 191426 444894
rect 191662 444658 227426 444894
rect 227662 444658 263426 444894
rect 263662 444658 299426 444894
rect 299662 444658 335426 444894
rect 335662 444658 371426 444894
rect 371662 444658 407426 444894
rect 407662 444658 443426 444894
rect 443662 444658 479426 444894
rect 479662 444658 515426 444894
rect 515662 444658 551426 444894
rect 551662 444658 591022 444894
rect 591258 444658 592350 444894
rect -8426 444574 592350 444658
rect -8426 444338 -7334 444574
rect -7098 444338 11426 444574
rect 11662 444338 47426 444574
rect 47662 444338 83426 444574
rect 83662 444338 119426 444574
rect 119662 444338 155426 444574
rect 155662 444338 191426 444574
rect 191662 444338 227426 444574
rect 227662 444338 263426 444574
rect 263662 444338 299426 444574
rect 299662 444338 335426 444574
rect 335662 444338 371426 444574
rect 371662 444338 407426 444574
rect 407662 444338 443426 444574
rect 443662 444338 479426 444574
rect 479662 444338 515426 444574
rect 515662 444338 551426 444574
rect 551662 444338 591022 444574
rect 591258 444338 592350 444574
rect -8426 444326 592350 444338
rect -7506 444314 -6926 444326
rect 11254 444314 11834 444326
rect 47254 444314 47834 444326
rect 83254 444314 83834 444326
rect 119254 444314 119834 444326
rect 155254 444314 155834 444326
rect 191254 444314 191834 444326
rect 227254 444314 227834 444326
rect 263254 444314 263834 444326
rect 299254 444314 299834 444326
rect 335254 444314 335834 444326
rect 371254 444314 371834 444326
rect 407254 444314 407834 444326
rect 443254 444314 443834 444326
rect 479254 444314 479834 444326
rect 515254 444314 515834 444326
rect 551254 444314 551834 444326
rect 590850 444314 591430 444326
rect -5666 441426 -5086 441438
rect 7774 441426 8354 441438
rect 43774 441426 44354 441438
rect 79774 441426 80354 441438
rect 115774 441426 116354 441438
rect 151774 441426 152354 441438
rect 187774 441426 188354 441438
rect 223774 441426 224354 441438
rect 259774 441426 260354 441438
rect 295774 441426 296354 441438
rect 331774 441426 332354 441438
rect 367774 441426 368354 441438
rect 403774 441426 404354 441438
rect 439774 441426 440354 441438
rect 475774 441426 476354 441438
rect 511774 441426 512354 441438
rect 547774 441426 548354 441438
rect 589010 441426 589590 441438
rect -6586 441414 590510 441426
rect -6586 441178 -5494 441414
rect -5258 441178 7946 441414
rect 8182 441178 43946 441414
rect 44182 441178 79946 441414
rect 80182 441178 115946 441414
rect 116182 441178 151946 441414
rect 152182 441178 187946 441414
rect 188182 441178 223946 441414
rect 224182 441178 259946 441414
rect 260182 441178 295946 441414
rect 296182 441178 331946 441414
rect 332182 441178 367946 441414
rect 368182 441178 403946 441414
rect 404182 441178 439946 441414
rect 440182 441178 475946 441414
rect 476182 441178 511946 441414
rect 512182 441178 547946 441414
rect 548182 441178 589182 441414
rect 589418 441178 590510 441414
rect -6586 441094 590510 441178
rect -6586 440858 -5494 441094
rect -5258 440858 7946 441094
rect 8182 440858 43946 441094
rect 44182 440858 79946 441094
rect 80182 440858 115946 441094
rect 116182 440858 151946 441094
rect 152182 440858 187946 441094
rect 188182 440858 223946 441094
rect 224182 440858 259946 441094
rect 260182 440858 295946 441094
rect 296182 440858 331946 441094
rect 332182 440858 367946 441094
rect 368182 440858 403946 441094
rect 404182 440858 439946 441094
rect 440182 440858 475946 441094
rect 476182 440858 511946 441094
rect 512182 440858 547946 441094
rect 548182 440858 589182 441094
rect 589418 440858 590510 441094
rect -6586 440846 590510 440858
rect -5666 440834 -5086 440846
rect 7774 440834 8354 440846
rect 43774 440834 44354 440846
rect 79774 440834 80354 440846
rect 115774 440834 116354 440846
rect 151774 440834 152354 440846
rect 187774 440834 188354 440846
rect 223774 440834 224354 440846
rect 259774 440834 260354 440846
rect 295774 440834 296354 440846
rect 331774 440834 332354 440846
rect 367774 440834 368354 440846
rect 403774 440834 404354 440846
rect 439774 440834 440354 440846
rect 475774 440834 476354 440846
rect 511774 440834 512354 440846
rect 547774 440834 548354 440846
rect 589010 440834 589590 440846
rect -3826 437946 -3246 437958
rect 4294 437946 4874 437958
rect 40294 437946 40874 437958
rect 76294 437946 76874 437958
rect 112294 437946 112874 437958
rect 148294 437946 148874 437958
rect 184294 437946 184874 437958
rect 220294 437946 220874 437958
rect 256294 437946 256874 437958
rect 292294 437946 292874 437958
rect 328294 437946 328874 437958
rect 364294 437946 364874 437958
rect 400294 437946 400874 437958
rect 436294 437946 436874 437958
rect 472294 437946 472874 437958
rect 508294 437946 508874 437958
rect 544294 437946 544874 437958
rect 580294 437946 580874 437958
rect 587170 437946 587750 437958
rect -4746 437934 588670 437946
rect -4746 437698 -3654 437934
rect -3418 437698 4466 437934
rect 4702 437698 40466 437934
rect 40702 437698 76466 437934
rect 76702 437698 112466 437934
rect 112702 437698 148466 437934
rect 148702 437698 184466 437934
rect 184702 437698 220466 437934
rect 220702 437698 256466 437934
rect 256702 437698 292466 437934
rect 292702 437698 328466 437934
rect 328702 437698 364466 437934
rect 364702 437698 400466 437934
rect 400702 437698 436466 437934
rect 436702 437698 472466 437934
rect 472702 437698 508466 437934
rect 508702 437698 544466 437934
rect 544702 437698 580466 437934
rect 580702 437698 587342 437934
rect 587578 437698 588670 437934
rect -4746 437614 588670 437698
rect -4746 437378 -3654 437614
rect -3418 437378 4466 437614
rect 4702 437378 40466 437614
rect 40702 437378 76466 437614
rect 76702 437378 112466 437614
rect 112702 437378 148466 437614
rect 148702 437378 184466 437614
rect 184702 437378 220466 437614
rect 220702 437378 256466 437614
rect 256702 437378 292466 437614
rect 292702 437378 328466 437614
rect 328702 437378 364466 437614
rect 364702 437378 400466 437614
rect 400702 437378 436466 437614
rect 436702 437378 472466 437614
rect 472702 437378 508466 437614
rect 508702 437378 544466 437614
rect 544702 437378 580466 437614
rect 580702 437378 587342 437614
rect 587578 437378 588670 437614
rect -4746 437366 588670 437378
rect -3826 437354 -3246 437366
rect 4294 437354 4874 437366
rect 40294 437354 40874 437366
rect 76294 437354 76874 437366
rect 112294 437354 112874 437366
rect 148294 437354 148874 437366
rect 184294 437354 184874 437366
rect 220294 437354 220874 437366
rect 256294 437354 256874 437366
rect 292294 437354 292874 437366
rect 328294 437354 328874 437366
rect 364294 437354 364874 437366
rect 400294 437354 400874 437366
rect 436294 437354 436874 437366
rect 472294 437354 472874 437366
rect 508294 437354 508874 437366
rect 544294 437354 544874 437366
rect 580294 437354 580874 437366
rect 587170 437354 587750 437366
rect -1986 434466 -1406 434478
rect 814 434466 1394 434478
rect 36814 434466 37394 434478
rect 72814 434466 73394 434478
rect 108814 434466 109394 434478
rect 144814 434466 145394 434478
rect 180814 434466 181394 434478
rect 216814 434466 217394 434478
rect 252814 434466 253394 434478
rect 288814 434466 289394 434478
rect 324814 434466 325394 434478
rect 360814 434466 361394 434478
rect 396814 434466 397394 434478
rect 432814 434466 433394 434478
rect 468814 434466 469394 434478
rect 504814 434466 505394 434478
rect 540814 434466 541394 434478
rect 576814 434466 577394 434478
rect 585330 434466 585910 434478
rect -2906 434454 586830 434466
rect -2906 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586830 434454
rect -2906 434134 586830 434218
rect -2906 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586830 434134
rect -2906 433886 586830 433898
rect -1986 433874 -1406 433886
rect 814 433874 1394 433886
rect 36814 433874 37394 433886
rect 72814 433874 73394 433886
rect 108814 433874 109394 433886
rect 144814 433874 145394 433886
rect 180814 433874 181394 433886
rect 216814 433874 217394 433886
rect 252814 433874 253394 433886
rect 288814 433874 289394 433886
rect 324814 433874 325394 433886
rect 360814 433874 361394 433886
rect 396814 433874 397394 433886
rect 432814 433874 433394 433886
rect 468814 433874 469394 433886
rect 504814 433874 505394 433886
rect 540814 433874 541394 433886
rect 576814 433874 577394 433886
rect 585330 433874 585910 433886
rect -8426 426906 -7846 426918
rect 29254 426906 29834 426918
rect 65254 426906 65834 426918
rect 101254 426906 101834 426918
rect 137254 426906 137834 426918
rect 173254 426906 173834 426918
rect 209254 426906 209834 426918
rect 245254 426906 245834 426918
rect 281254 426906 281834 426918
rect 317254 426906 317834 426918
rect 353254 426906 353834 426918
rect 389254 426906 389834 426918
rect 425254 426906 425834 426918
rect 461254 426906 461834 426918
rect 497254 426906 497834 426918
rect 533254 426906 533834 426918
rect 569254 426906 569834 426918
rect 591770 426906 592350 426918
rect -8426 426894 592350 426906
rect -8426 426658 -8254 426894
rect -8018 426658 29426 426894
rect 29662 426658 65426 426894
rect 65662 426658 101426 426894
rect 101662 426658 137426 426894
rect 137662 426658 173426 426894
rect 173662 426658 209426 426894
rect 209662 426658 245426 426894
rect 245662 426658 281426 426894
rect 281662 426658 317426 426894
rect 317662 426658 353426 426894
rect 353662 426658 389426 426894
rect 389662 426658 425426 426894
rect 425662 426658 461426 426894
rect 461662 426658 497426 426894
rect 497662 426658 533426 426894
rect 533662 426658 569426 426894
rect 569662 426658 591942 426894
rect 592178 426658 592350 426894
rect -8426 426574 592350 426658
rect -8426 426338 -8254 426574
rect -8018 426338 29426 426574
rect 29662 426338 65426 426574
rect 65662 426338 101426 426574
rect 101662 426338 137426 426574
rect 137662 426338 173426 426574
rect 173662 426338 209426 426574
rect 209662 426338 245426 426574
rect 245662 426338 281426 426574
rect 281662 426338 317426 426574
rect 317662 426338 353426 426574
rect 353662 426338 389426 426574
rect 389662 426338 425426 426574
rect 425662 426338 461426 426574
rect 461662 426338 497426 426574
rect 497662 426338 533426 426574
rect 533662 426338 569426 426574
rect 569662 426338 591942 426574
rect 592178 426338 592350 426574
rect -8426 426326 592350 426338
rect -8426 426314 -7846 426326
rect 29254 426314 29834 426326
rect 65254 426314 65834 426326
rect 101254 426314 101834 426326
rect 137254 426314 137834 426326
rect 173254 426314 173834 426326
rect 209254 426314 209834 426326
rect 245254 426314 245834 426326
rect 281254 426314 281834 426326
rect 317254 426314 317834 426326
rect 353254 426314 353834 426326
rect 389254 426314 389834 426326
rect 425254 426314 425834 426326
rect 461254 426314 461834 426326
rect 497254 426314 497834 426326
rect 533254 426314 533834 426326
rect 569254 426314 569834 426326
rect 591770 426314 592350 426326
rect -6586 423426 -6006 423438
rect 25774 423426 26354 423438
rect 61774 423426 62354 423438
rect 97774 423426 98354 423438
rect 133774 423426 134354 423438
rect 169774 423426 170354 423438
rect 205774 423426 206354 423438
rect 241774 423426 242354 423438
rect 277774 423426 278354 423438
rect 313774 423426 314354 423438
rect 349774 423426 350354 423438
rect 385774 423426 386354 423438
rect 421774 423426 422354 423438
rect 457774 423426 458354 423438
rect 493774 423426 494354 423438
rect 529774 423426 530354 423438
rect 565774 423426 566354 423438
rect 589930 423426 590510 423438
rect -6586 423414 590510 423426
rect -6586 423178 -6414 423414
rect -6178 423178 25946 423414
rect 26182 423178 61946 423414
rect 62182 423178 97946 423414
rect 98182 423178 133946 423414
rect 134182 423178 169946 423414
rect 170182 423178 205946 423414
rect 206182 423178 241946 423414
rect 242182 423178 277946 423414
rect 278182 423178 313946 423414
rect 314182 423178 349946 423414
rect 350182 423178 385946 423414
rect 386182 423178 421946 423414
rect 422182 423178 457946 423414
rect 458182 423178 493946 423414
rect 494182 423178 529946 423414
rect 530182 423178 565946 423414
rect 566182 423178 590102 423414
rect 590338 423178 590510 423414
rect -6586 423094 590510 423178
rect -6586 422858 -6414 423094
rect -6178 422858 25946 423094
rect 26182 422858 61946 423094
rect 62182 422858 97946 423094
rect 98182 422858 133946 423094
rect 134182 422858 169946 423094
rect 170182 422858 205946 423094
rect 206182 422858 241946 423094
rect 242182 422858 277946 423094
rect 278182 422858 313946 423094
rect 314182 422858 349946 423094
rect 350182 422858 385946 423094
rect 386182 422858 421946 423094
rect 422182 422858 457946 423094
rect 458182 422858 493946 423094
rect 494182 422858 529946 423094
rect 530182 422858 565946 423094
rect 566182 422858 590102 423094
rect 590338 422858 590510 423094
rect -6586 422846 590510 422858
rect -6586 422834 -6006 422846
rect 25774 422834 26354 422846
rect 61774 422834 62354 422846
rect 97774 422834 98354 422846
rect 133774 422834 134354 422846
rect 169774 422834 170354 422846
rect 205774 422834 206354 422846
rect 241774 422834 242354 422846
rect 277774 422834 278354 422846
rect 313774 422834 314354 422846
rect 349774 422834 350354 422846
rect 385774 422834 386354 422846
rect 421774 422834 422354 422846
rect 457774 422834 458354 422846
rect 493774 422834 494354 422846
rect 529774 422834 530354 422846
rect 565774 422834 566354 422846
rect 589930 422834 590510 422846
rect -4746 419946 -4166 419958
rect 22294 419946 22874 419958
rect 58294 419946 58874 419958
rect 94294 419946 94874 419958
rect 130294 419946 130874 419958
rect 166294 419946 166874 419958
rect 202294 419946 202874 419958
rect 238294 419946 238874 419958
rect 274294 419946 274874 419958
rect 310294 419946 310874 419958
rect 346294 419946 346874 419958
rect 382294 419946 382874 419958
rect 418294 419946 418874 419958
rect 454294 419946 454874 419958
rect 490294 419946 490874 419958
rect 526294 419946 526874 419958
rect 562294 419946 562874 419958
rect 588090 419946 588670 419958
rect -4746 419934 588670 419946
rect -4746 419698 -4574 419934
rect -4338 419698 22466 419934
rect 22702 419698 58466 419934
rect 58702 419698 94466 419934
rect 94702 419698 130466 419934
rect 130702 419698 166466 419934
rect 166702 419698 202466 419934
rect 202702 419698 238466 419934
rect 238702 419698 274466 419934
rect 274702 419698 310466 419934
rect 310702 419698 346466 419934
rect 346702 419698 382466 419934
rect 382702 419698 418466 419934
rect 418702 419698 454466 419934
rect 454702 419698 490466 419934
rect 490702 419698 526466 419934
rect 526702 419698 562466 419934
rect 562702 419698 588262 419934
rect 588498 419698 588670 419934
rect -4746 419614 588670 419698
rect -4746 419378 -4574 419614
rect -4338 419378 22466 419614
rect 22702 419378 58466 419614
rect 58702 419378 94466 419614
rect 94702 419378 130466 419614
rect 130702 419378 166466 419614
rect 166702 419378 202466 419614
rect 202702 419378 238466 419614
rect 238702 419378 274466 419614
rect 274702 419378 310466 419614
rect 310702 419378 346466 419614
rect 346702 419378 382466 419614
rect 382702 419378 418466 419614
rect 418702 419378 454466 419614
rect 454702 419378 490466 419614
rect 490702 419378 526466 419614
rect 526702 419378 562466 419614
rect 562702 419378 588262 419614
rect 588498 419378 588670 419614
rect -4746 419366 588670 419378
rect -4746 419354 -4166 419366
rect 22294 419354 22874 419366
rect 58294 419354 58874 419366
rect 94294 419354 94874 419366
rect 130294 419354 130874 419366
rect 166294 419354 166874 419366
rect 202294 419354 202874 419366
rect 238294 419354 238874 419366
rect 274294 419354 274874 419366
rect 310294 419354 310874 419366
rect 346294 419354 346874 419366
rect 382294 419354 382874 419366
rect 418294 419354 418874 419366
rect 454294 419354 454874 419366
rect 490294 419354 490874 419366
rect 526294 419354 526874 419366
rect 562294 419354 562874 419366
rect 588090 419354 588670 419366
rect -2906 416466 -2326 416478
rect 18814 416466 19394 416478
rect 54814 416466 55394 416478
rect 90814 416466 91394 416478
rect 126814 416466 127394 416478
rect 162814 416466 163394 416478
rect 198814 416466 199394 416478
rect 234814 416466 235394 416478
rect 270814 416466 271394 416478
rect 306814 416466 307394 416478
rect 342814 416466 343394 416478
rect 378814 416466 379394 416478
rect 414814 416466 415394 416478
rect 450814 416466 451394 416478
rect 486814 416466 487394 416478
rect 522814 416466 523394 416478
rect 558814 416466 559394 416478
rect 586250 416466 586830 416478
rect -2906 416454 586830 416466
rect -2906 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586830 416454
rect -2906 416134 586830 416218
rect -2906 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586830 416134
rect -2906 415886 586830 415898
rect -2906 415874 -2326 415886
rect 18814 415874 19394 415886
rect 54814 415874 55394 415886
rect 90814 415874 91394 415886
rect 126814 415874 127394 415886
rect 162814 415874 163394 415886
rect 198814 415874 199394 415886
rect 234814 415874 235394 415886
rect 270814 415874 271394 415886
rect 306814 415874 307394 415886
rect 342814 415874 343394 415886
rect 378814 415874 379394 415886
rect 414814 415874 415394 415886
rect 450814 415874 451394 415886
rect 486814 415874 487394 415886
rect 522814 415874 523394 415886
rect 558814 415874 559394 415886
rect 586250 415874 586830 415886
rect -7506 408906 -6926 408918
rect 11254 408906 11834 408918
rect 47254 408906 47834 408918
rect 83254 408906 83834 408918
rect 119254 408906 119834 408918
rect 155254 408906 155834 408918
rect 191254 408906 191834 408918
rect 227254 408906 227834 408918
rect 263254 408906 263834 408918
rect 299254 408906 299834 408918
rect 335254 408906 335834 408918
rect 371254 408906 371834 408918
rect 407254 408906 407834 408918
rect 443254 408906 443834 408918
rect 479254 408906 479834 408918
rect 515254 408906 515834 408918
rect 551254 408906 551834 408918
rect 590850 408906 591430 408918
rect -8426 408894 592350 408906
rect -8426 408658 -7334 408894
rect -7098 408658 11426 408894
rect 11662 408658 47426 408894
rect 47662 408658 83426 408894
rect 83662 408658 119426 408894
rect 119662 408658 155426 408894
rect 155662 408658 191426 408894
rect 191662 408658 227426 408894
rect 227662 408658 263426 408894
rect 263662 408658 299426 408894
rect 299662 408658 335426 408894
rect 335662 408658 371426 408894
rect 371662 408658 407426 408894
rect 407662 408658 443426 408894
rect 443662 408658 479426 408894
rect 479662 408658 515426 408894
rect 515662 408658 551426 408894
rect 551662 408658 591022 408894
rect 591258 408658 592350 408894
rect -8426 408574 592350 408658
rect -8426 408338 -7334 408574
rect -7098 408338 11426 408574
rect 11662 408338 47426 408574
rect 47662 408338 83426 408574
rect 83662 408338 119426 408574
rect 119662 408338 155426 408574
rect 155662 408338 191426 408574
rect 191662 408338 227426 408574
rect 227662 408338 263426 408574
rect 263662 408338 299426 408574
rect 299662 408338 335426 408574
rect 335662 408338 371426 408574
rect 371662 408338 407426 408574
rect 407662 408338 443426 408574
rect 443662 408338 479426 408574
rect 479662 408338 515426 408574
rect 515662 408338 551426 408574
rect 551662 408338 591022 408574
rect 591258 408338 592350 408574
rect -8426 408326 592350 408338
rect -7506 408314 -6926 408326
rect 11254 408314 11834 408326
rect 47254 408314 47834 408326
rect 83254 408314 83834 408326
rect 119254 408314 119834 408326
rect 155254 408314 155834 408326
rect 191254 408314 191834 408326
rect 227254 408314 227834 408326
rect 263254 408314 263834 408326
rect 299254 408314 299834 408326
rect 335254 408314 335834 408326
rect 371254 408314 371834 408326
rect 407254 408314 407834 408326
rect 443254 408314 443834 408326
rect 479254 408314 479834 408326
rect 515254 408314 515834 408326
rect 551254 408314 551834 408326
rect 590850 408314 591430 408326
rect -5666 405426 -5086 405438
rect 7774 405426 8354 405438
rect 43774 405426 44354 405438
rect 79774 405426 80354 405438
rect 115774 405426 116354 405438
rect 151774 405426 152354 405438
rect 187774 405426 188354 405438
rect 223774 405426 224354 405438
rect 259774 405426 260354 405438
rect 295774 405426 296354 405438
rect 331774 405426 332354 405438
rect 367774 405426 368354 405438
rect 403774 405426 404354 405438
rect 439774 405426 440354 405438
rect 475774 405426 476354 405438
rect 511774 405426 512354 405438
rect 547774 405426 548354 405438
rect 589010 405426 589590 405438
rect -6586 405414 590510 405426
rect -6586 405178 -5494 405414
rect -5258 405178 7946 405414
rect 8182 405178 43946 405414
rect 44182 405178 79946 405414
rect 80182 405178 115946 405414
rect 116182 405178 151946 405414
rect 152182 405178 187946 405414
rect 188182 405178 223946 405414
rect 224182 405178 259946 405414
rect 260182 405178 295946 405414
rect 296182 405178 331946 405414
rect 332182 405178 367946 405414
rect 368182 405178 403946 405414
rect 404182 405178 439946 405414
rect 440182 405178 475946 405414
rect 476182 405178 511946 405414
rect 512182 405178 547946 405414
rect 548182 405178 589182 405414
rect 589418 405178 590510 405414
rect -6586 405094 590510 405178
rect -6586 404858 -5494 405094
rect -5258 404858 7946 405094
rect 8182 404858 43946 405094
rect 44182 404858 79946 405094
rect 80182 404858 115946 405094
rect 116182 404858 151946 405094
rect 152182 404858 187946 405094
rect 188182 404858 223946 405094
rect 224182 404858 259946 405094
rect 260182 404858 295946 405094
rect 296182 404858 331946 405094
rect 332182 404858 367946 405094
rect 368182 404858 403946 405094
rect 404182 404858 439946 405094
rect 440182 404858 475946 405094
rect 476182 404858 511946 405094
rect 512182 404858 547946 405094
rect 548182 404858 589182 405094
rect 589418 404858 590510 405094
rect -6586 404846 590510 404858
rect -5666 404834 -5086 404846
rect 7774 404834 8354 404846
rect 43774 404834 44354 404846
rect 79774 404834 80354 404846
rect 115774 404834 116354 404846
rect 151774 404834 152354 404846
rect 187774 404834 188354 404846
rect 223774 404834 224354 404846
rect 259774 404834 260354 404846
rect 295774 404834 296354 404846
rect 331774 404834 332354 404846
rect 367774 404834 368354 404846
rect 403774 404834 404354 404846
rect 439774 404834 440354 404846
rect 475774 404834 476354 404846
rect 511774 404834 512354 404846
rect 547774 404834 548354 404846
rect 589010 404834 589590 404846
rect -3826 401946 -3246 401958
rect 4294 401946 4874 401958
rect 40294 401946 40874 401958
rect 76294 401946 76874 401958
rect 112294 401946 112874 401958
rect 148294 401946 148874 401958
rect 184294 401946 184874 401958
rect 220294 401946 220874 401958
rect 256294 401946 256874 401958
rect 292294 401946 292874 401958
rect 328294 401946 328874 401958
rect 364294 401946 364874 401958
rect 400294 401946 400874 401958
rect 436294 401946 436874 401958
rect 472294 401946 472874 401958
rect 508294 401946 508874 401958
rect 544294 401946 544874 401958
rect 580294 401946 580874 401958
rect 587170 401946 587750 401958
rect -4746 401934 588670 401946
rect -4746 401698 -3654 401934
rect -3418 401698 4466 401934
rect 4702 401698 40466 401934
rect 40702 401698 76466 401934
rect 76702 401698 112466 401934
rect 112702 401698 148466 401934
rect 148702 401698 184466 401934
rect 184702 401698 220466 401934
rect 220702 401698 256466 401934
rect 256702 401698 292466 401934
rect 292702 401698 328466 401934
rect 328702 401698 364466 401934
rect 364702 401698 400466 401934
rect 400702 401698 436466 401934
rect 436702 401698 472466 401934
rect 472702 401698 508466 401934
rect 508702 401698 544466 401934
rect 544702 401698 580466 401934
rect 580702 401698 587342 401934
rect 587578 401698 588670 401934
rect -4746 401614 588670 401698
rect -4746 401378 -3654 401614
rect -3418 401378 4466 401614
rect 4702 401378 40466 401614
rect 40702 401378 76466 401614
rect 76702 401378 112466 401614
rect 112702 401378 148466 401614
rect 148702 401378 184466 401614
rect 184702 401378 220466 401614
rect 220702 401378 256466 401614
rect 256702 401378 292466 401614
rect 292702 401378 328466 401614
rect 328702 401378 364466 401614
rect 364702 401378 400466 401614
rect 400702 401378 436466 401614
rect 436702 401378 472466 401614
rect 472702 401378 508466 401614
rect 508702 401378 544466 401614
rect 544702 401378 580466 401614
rect 580702 401378 587342 401614
rect 587578 401378 588670 401614
rect -4746 401366 588670 401378
rect -3826 401354 -3246 401366
rect 4294 401354 4874 401366
rect 40294 401354 40874 401366
rect 76294 401354 76874 401366
rect 112294 401354 112874 401366
rect 148294 401354 148874 401366
rect 184294 401354 184874 401366
rect 220294 401354 220874 401366
rect 256294 401354 256874 401366
rect 292294 401354 292874 401366
rect 328294 401354 328874 401366
rect 364294 401354 364874 401366
rect 400294 401354 400874 401366
rect 436294 401354 436874 401366
rect 472294 401354 472874 401366
rect 508294 401354 508874 401366
rect 544294 401354 544874 401366
rect 580294 401354 580874 401366
rect 587170 401354 587750 401366
rect -1986 398466 -1406 398478
rect 814 398466 1394 398478
rect 36814 398466 37394 398478
rect 72814 398466 73394 398478
rect 108814 398466 109394 398478
rect 144814 398466 145394 398478
rect 180814 398466 181394 398478
rect 216814 398466 217394 398478
rect 252814 398466 253394 398478
rect 288814 398466 289394 398478
rect 324814 398466 325394 398478
rect 360814 398466 361394 398478
rect 396814 398466 397394 398478
rect 432814 398466 433394 398478
rect 468814 398466 469394 398478
rect 504814 398466 505394 398478
rect 540814 398466 541394 398478
rect 576814 398466 577394 398478
rect 585330 398466 585910 398478
rect -2906 398454 586830 398466
rect -2906 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586830 398454
rect -2906 398134 586830 398218
rect -2906 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586830 398134
rect -2906 397886 586830 397898
rect -1986 397874 -1406 397886
rect 814 397874 1394 397886
rect 36814 397874 37394 397886
rect 72814 397874 73394 397886
rect 108814 397874 109394 397886
rect 144814 397874 145394 397886
rect 180814 397874 181394 397886
rect 216814 397874 217394 397886
rect 252814 397874 253394 397886
rect 288814 397874 289394 397886
rect 324814 397874 325394 397886
rect 360814 397874 361394 397886
rect 396814 397874 397394 397886
rect 432814 397874 433394 397886
rect 468814 397874 469394 397886
rect 504814 397874 505394 397886
rect 540814 397874 541394 397886
rect 576814 397874 577394 397886
rect 585330 397874 585910 397886
rect -8426 390906 -7846 390918
rect 29254 390906 29834 390918
rect 65254 390906 65834 390918
rect 101254 390906 101834 390918
rect 137254 390906 137834 390918
rect 173254 390906 173834 390918
rect 209254 390906 209834 390918
rect 245254 390906 245834 390918
rect 281254 390906 281834 390918
rect 317254 390906 317834 390918
rect 353254 390906 353834 390918
rect 389254 390906 389834 390918
rect 425254 390906 425834 390918
rect 461254 390906 461834 390918
rect 497254 390906 497834 390918
rect 533254 390906 533834 390918
rect 569254 390906 569834 390918
rect 591770 390906 592350 390918
rect -8426 390894 592350 390906
rect -8426 390658 -8254 390894
rect -8018 390658 29426 390894
rect 29662 390658 65426 390894
rect 65662 390658 101426 390894
rect 101662 390658 137426 390894
rect 137662 390658 173426 390894
rect 173662 390658 209426 390894
rect 209662 390658 245426 390894
rect 245662 390658 281426 390894
rect 281662 390658 317426 390894
rect 317662 390658 353426 390894
rect 353662 390658 389426 390894
rect 389662 390658 425426 390894
rect 425662 390658 461426 390894
rect 461662 390658 497426 390894
rect 497662 390658 533426 390894
rect 533662 390658 569426 390894
rect 569662 390658 591942 390894
rect 592178 390658 592350 390894
rect -8426 390574 592350 390658
rect -8426 390338 -8254 390574
rect -8018 390338 29426 390574
rect 29662 390338 65426 390574
rect 65662 390338 101426 390574
rect 101662 390338 137426 390574
rect 137662 390338 173426 390574
rect 173662 390338 209426 390574
rect 209662 390338 245426 390574
rect 245662 390338 281426 390574
rect 281662 390338 317426 390574
rect 317662 390338 353426 390574
rect 353662 390338 389426 390574
rect 389662 390338 425426 390574
rect 425662 390338 461426 390574
rect 461662 390338 497426 390574
rect 497662 390338 533426 390574
rect 533662 390338 569426 390574
rect 569662 390338 591942 390574
rect 592178 390338 592350 390574
rect -8426 390326 592350 390338
rect -8426 390314 -7846 390326
rect 29254 390314 29834 390326
rect 65254 390314 65834 390326
rect 101254 390314 101834 390326
rect 137254 390314 137834 390326
rect 173254 390314 173834 390326
rect 209254 390314 209834 390326
rect 245254 390314 245834 390326
rect 281254 390314 281834 390326
rect 317254 390314 317834 390326
rect 353254 390314 353834 390326
rect 389254 390314 389834 390326
rect 425254 390314 425834 390326
rect 461254 390314 461834 390326
rect 497254 390314 497834 390326
rect 533254 390314 533834 390326
rect 569254 390314 569834 390326
rect 591770 390314 592350 390326
rect -6586 387426 -6006 387438
rect 25774 387426 26354 387438
rect 61774 387426 62354 387438
rect 97774 387426 98354 387438
rect 133774 387426 134354 387438
rect 169774 387426 170354 387438
rect 205774 387426 206354 387438
rect 241774 387426 242354 387438
rect 277774 387426 278354 387438
rect 313774 387426 314354 387438
rect 349774 387426 350354 387438
rect 385774 387426 386354 387438
rect 421774 387426 422354 387438
rect 457774 387426 458354 387438
rect 493774 387426 494354 387438
rect 529774 387426 530354 387438
rect 565774 387426 566354 387438
rect 589930 387426 590510 387438
rect -6586 387414 590510 387426
rect -6586 387178 -6414 387414
rect -6178 387178 25946 387414
rect 26182 387178 61946 387414
rect 62182 387178 97946 387414
rect 98182 387178 133946 387414
rect 134182 387178 169946 387414
rect 170182 387178 205946 387414
rect 206182 387178 241946 387414
rect 242182 387178 277946 387414
rect 278182 387178 313946 387414
rect 314182 387178 349946 387414
rect 350182 387178 385946 387414
rect 386182 387178 421946 387414
rect 422182 387178 457946 387414
rect 458182 387178 493946 387414
rect 494182 387178 529946 387414
rect 530182 387178 565946 387414
rect 566182 387178 590102 387414
rect 590338 387178 590510 387414
rect -6586 387094 590510 387178
rect -6586 386858 -6414 387094
rect -6178 386858 25946 387094
rect 26182 386858 61946 387094
rect 62182 386858 97946 387094
rect 98182 386858 133946 387094
rect 134182 386858 169946 387094
rect 170182 386858 205946 387094
rect 206182 386858 241946 387094
rect 242182 386858 277946 387094
rect 278182 386858 313946 387094
rect 314182 386858 349946 387094
rect 350182 386858 385946 387094
rect 386182 386858 421946 387094
rect 422182 386858 457946 387094
rect 458182 386858 493946 387094
rect 494182 386858 529946 387094
rect 530182 386858 565946 387094
rect 566182 386858 590102 387094
rect 590338 386858 590510 387094
rect -6586 386846 590510 386858
rect -6586 386834 -6006 386846
rect 25774 386834 26354 386846
rect 61774 386834 62354 386846
rect 97774 386834 98354 386846
rect 133774 386834 134354 386846
rect 169774 386834 170354 386846
rect 205774 386834 206354 386846
rect 241774 386834 242354 386846
rect 277774 386834 278354 386846
rect 313774 386834 314354 386846
rect 349774 386834 350354 386846
rect 385774 386834 386354 386846
rect 421774 386834 422354 386846
rect 457774 386834 458354 386846
rect 493774 386834 494354 386846
rect 529774 386834 530354 386846
rect 565774 386834 566354 386846
rect 589930 386834 590510 386846
rect -4746 383946 -4166 383958
rect 22294 383946 22874 383958
rect 58294 383946 58874 383958
rect 94294 383946 94874 383958
rect 130294 383946 130874 383958
rect 166294 383946 166874 383958
rect 202294 383946 202874 383958
rect 238294 383946 238874 383958
rect 274294 383946 274874 383958
rect 310294 383946 310874 383958
rect 346294 383946 346874 383958
rect 382294 383946 382874 383958
rect 418294 383946 418874 383958
rect 454294 383946 454874 383958
rect 490294 383946 490874 383958
rect 526294 383946 526874 383958
rect 562294 383946 562874 383958
rect 588090 383946 588670 383958
rect -4746 383934 588670 383946
rect -4746 383698 -4574 383934
rect -4338 383698 22466 383934
rect 22702 383698 58466 383934
rect 58702 383698 94466 383934
rect 94702 383698 130466 383934
rect 130702 383698 166466 383934
rect 166702 383698 202466 383934
rect 202702 383698 238466 383934
rect 238702 383698 274466 383934
rect 274702 383698 310466 383934
rect 310702 383698 346466 383934
rect 346702 383698 382466 383934
rect 382702 383698 418466 383934
rect 418702 383698 454466 383934
rect 454702 383698 490466 383934
rect 490702 383698 526466 383934
rect 526702 383698 562466 383934
rect 562702 383698 588262 383934
rect 588498 383698 588670 383934
rect -4746 383614 588670 383698
rect -4746 383378 -4574 383614
rect -4338 383378 22466 383614
rect 22702 383378 58466 383614
rect 58702 383378 94466 383614
rect 94702 383378 130466 383614
rect 130702 383378 166466 383614
rect 166702 383378 202466 383614
rect 202702 383378 238466 383614
rect 238702 383378 274466 383614
rect 274702 383378 310466 383614
rect 310702 383378 346466 383614
rect 346702 383378 382466 383614
rect 382702 383378 418466 383614
rect 418702 383378 454466 383614
rect 454702 383378 490466 383614
rect 490702 383378 526466 383614
rect 526702 383378 562466 383614
rect 562702 383378 588262 383614
rect 588498 383378 588670 383614
rect -4746 383366 588670 383378
rect -4746 383354 -4166 383366
rect 22294 383354 22874 383366
rect 58294 383354 58874 383366
rect 94294 383354 94874 383366
rect 130294 383354 130874 383366
rect 166294 383354 166874 383366
rect 202294 383354 202874 383366
rect 238294 383354 238874 383366
rect 274294 383354 274874 383366
rect 310294 383354 310874 383366
rect 346294 383354 346874 383366
rect 382294 383354 382874 383366
rect 418294 383354 418874 383366
rect 454294 383354 454874 383366
rect 490294 383354 490874 383366
rect 526294 383354 526874 383366
rect 562294 383354 562874 383366
rect 588090 383354 588670 383366
rect -2906 380466 -2326 380478
rect 18814 380466 19394 380478
rect 54814 380466 55394 380478
rect 90814 380466 91394 380478
rect 126814 380466 127394 380478
rect 162814 380466 163394 380478
rect 198814 380466 199394 380478
rect 234814 380466 235394 380478
rect 270814 380466 271394 380478
rect 306814 380466 307394 380478
rect 342814 380466 343394 380478
rect 378814 380466 379394 380478
rect 414814 380466 415394 380478
rect 450814 380466 451394 380478
rect 486814 380466 487394 380478
rect 522814 380466 523394 380478
rect 558814 380466 559394 380478
rect 586250 380466 586830 380478
rect -2906 380454 586830 380466
rect -2906 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586830 380454
rect -2906 380134 586830 380218
rect -2906 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586830 380134
rect -2906 379886 586830 379898
rect -2906 379874 -2326 379886
rect 18814 379874 19394 379886
rect 54814 379874 55394 379886
rect 90814 379874 91394 379886
rect 126814 379874 127394 379886
rect 162814 379874 163394 379886
rect 198814 379874 199394 379886
rect 234814 379874 235394 379886
rect 270814 379874 271394 379886
rect 306814 379874 307394 379886
rect 342814 379874 343394 379886
rect 378814 379874 379394 379886
rect 414814 379874 415394 379886
rect 450814 379874 451394 379886
rect 486814 379874 487394 379886
rect 522814 379874 523394 379886
rect 558814 379874 559394 379886
rect 586250 379874 586830 379886
rect -7506 372906 -6926 372918
rect 11254 372906 11834 372918
rect 47254 372906 47834 372918
rect 83254 372906 83834 372918
rect 119254 372906 119834 372918
rect 155254 372906 155834 372918
rect 191254 372906 191834 372918
rect 227254 372906 227834 372918
rect 263254 372906 263834 372918
rect 299254 372906 299834 372918
rect 335254 372906 335834 372918
rect 371254 372906 371834 372918
rect 407254 372906 407834 372918
rect 443254 372906 443834 372918
rect 479254 372906 479834 372918
rect 515254 372906 515834 372918
rect 551254 372906 551834 372918
rect 590850 372906 591430 372918
rect -8426 372894 592350 372906
rect -8426 372658 -7334 372894
rect -7098 372658 11426 372894
rect 11662 372658 47426 372894
rect 47662 372658 83426 372894
rect 83662 372658 119426 372894
rect 119662 372658 155426 372894
rect 155662 372658 191426 372894
rect 191662 372658 227426 372894
rect 227662 372658 263426 372894
rect 263662 372658 299426 372894
rect 299662 372658 335426 372894
rect 335662 372658 371426 372894
rect 371662 372658 407426 372894
rect 407662 372658 443426 372894
rect 443662 372658 479426 372894
rect 479662 372658 515426 372894
rect 515662 372658 551426 372894
rect 551662 372658 591022 372894
rect 591258 372658 592350 372894
rect -8426 372574 592350 372658
rect -8426 372338 -7334 372574
rect -7098 372338 11426 372574
rect 11662 372338 47426 372574
rect 47662 372338 83426 372574
rect 83662 372338 119426 372574
rect 119662 372338 155426 372574
rect 155662 372338 191426 372574
rect 191662 372338 227426 372574
rect 227662 372338 263426 372574
rect 263662 372338 299426 372574
rect 299662 372338 335426 372574
rect 335662 372338 371426 372574
rect 371662 372338 407426 372574
rect 407662 372338 443426 372574
rect 443662 372338 479426 372574
rect 479662 372338 515426 372574
rect 515662 372338 551426 372574
rect 551662 372338 591022 372574
rect 591258 372338 592350 372574
rect -8426 372326 592350 372338
rect -7506 372314 -6926 372326
rect 11254 372314 11834 372326
rect 47254 372314 47834 372326
rect 83254 372314 83834 372326
rect 119254 372314 119834 372326
rect 155254 372314 155834 372326
rect 191254 372314 191834 372326
rect 227254 372314 227834 372326
rect 263254 372314 263834 372326
rect 299254 372314 299834 372326
rect 335254 372314 335834 372326
rect 371254 372314 371834 372326
rect 407254 372314 407834 372326
rect 443254 372314 443834 372326
rect 479254 372314 479834 372326
rect 515254 372314 515834 372326
rect 551254 372314 551834 372326
rect 590850 372314 591430 372326
rect -5666 369426 -5086 369438
rect 7774 369426 8354 369438
rect 43774 369426 44354 369438
rect 79774 369426 80354 369438
rect 115774 369426 116354 369438
rect 151774 369426 152354 369438
rect 187774 369426 188354 369438
rect 223774 369426 224354 369438
rect 259774 369426 260354 369438
rect 295774 369426 296354 369438
rect 331774 369426 332354 369438
rect 367774 369426 368354 369438
rect 403774 369426 404354 369438
rect 439774 369426 440354 369438
rect 475774 369426 476354 369438
rect 511774 369426 512354 369438
rect 547774 369426 548354 369438
rect 589010 369426 589590 369438
rect -6586 369414 590510 369426
rect -6586 369178 -5494 369414
rect -5258 369178 7946 369414
rect 8182 369178 43946 369414
rect 44182 369178 79946 369414
rect 80182 369178 115946 369414
rect 116182 369178 151946 369414
rect 152182 369178 187946 369414
rect 188182 369178 223946 369414
rect 224182 369178 259946 369414
rect 260182 369178 295946 369414
rect 296182 369178 331946 369414
rect 332182 369178 367946 369414
rect 368182 369178 403946 369414
rect 404182 369178 439946 369414
rect 440182 369178 475946 369414
rect 476182 369178 511946 369414
rect 512182 369178 547946 369414
rect 548182 369178 589182 369414
rect 589418 369178 590510 369414
rect -6586 369094 590510 369178
rect -6586 368858 -5494 369094
rect -5258 368858 7946 369094
rect 8182 368858 43946 369094
rect 44182 368858 79946 369094
rect 80182 368858 115946 369094
rect 116182 368858 151946 369094
rect 152182 368858 187946 369094
rect 188182 368858 223946 369094
rect 224182 368858 259946 369094
rect 260182 368858 295946 369094
rect 296182 368858 331946 369094
rect 332182 368858 367946 369094
rect 368182 368858 403946 369094
rect 404182 368858 439946 369094
rect 440182 368858 475946 369094
rect 476182 368858 511946 369094
rect 512182 368858 547946 369094
rect 548182 368858 589182 369094
rect 589418 368858 590510 369094
rect -6586 368846 590510 368858
rect -5666 368834 -5086 368846
rect 7774 368834 8354 368846
rect 43774 368834 44354 368846
rect 79774 368834 80354 368846
rect 115774 368834 116354 368846
rect 151774 368834 152354 368846
rect 187774 368834 188354 368846
rect 223774 368834 224354 368846
rect 259774 368834 260354 368846
rect 295774 368834 296354 368846
rect 331774 368834 332354 368846
rect 367774 368834 368354 368846
rect 403774 368834 404354 368846
rect 439774 368834 440354 368846
rect 475774 368834 476354 368846
rect 511774 368834 512354 368846
rect 547774 368834 548354 368846
rect 589010 368834 589590 368846
rect -3826 365946 -3246 365958
rect 4294 365946 4874 365958
rect 40294 365946 40874 365958
rect 76294 365946 76874 365958
rect 112294 365946 112874 365958
rect 148294 365946 148874 365958
rect 184294 365946 184874 365958
rect 220294 365946 220874 365958
rect 256294 365946 256874 365958
rect 292294 365946 292874 365958
rect 328294 365946 328874 365958
rect 364294 365946 364874 365958
rect 400294 365946 400874 365958
rect 436294 365946 436874 365958
rect 472294 365946 472874 365958
rect 508294 365946 508874 365958
rect 544294 365946 544874 365958
rect 580294 365946 580874 365958
rect 587170 365946 587750 365958
rect -4746 365934 588670 365946
rect -4746 365698 -3654 365934
rect -3418 365698 4466 365934
rect 4702 365698 40466 365934
rect 40702 365698 76466 365934
rect 76702 365698 112466 365934
rect 112702 365698 148466 365934
rect 148702 365698 184466 365934
rect 184702 365698 220466 365934
rect 220702 365698 256466 365934
rect 256702 365698 292466 365934
rect 292702 365698 328466 365934
rect 328702 365698 364466 365934
rect 364702 365698 400466 365934
rect 400702 365698 436466 365934
rect 436702 365698 472466 365934
rect 472702 365698 508466 365934
rect 508702 365698 544466 365934
rect 544702 365698 580466 365934
rect 580702 365698 587342 365934
rect 587578 365698 588670 365934
rect -4746 365614 588670 365698
rect -4746 365378 -3654 365614
rect -3418 365378 4466 365614
rect 4702 365378 40466 365614
rect 40702 365378 76466 365614
rect 76702 365378 112466 365614
rect 112702 365378 148466 365614
rect 148702 365378 184466 365614
rect 184702 365378 220466 365614
rect 220702 365378 256466 365614
rect 256702 365378 292466 365614
rect 292702 365378 328466 365614
rect 328702 365378 364466 365614
rect 364702 365378 400466 365614
rect 400702 365378 436466 365614
rect 436702 365378 472466 365614
rect 472702 365378 508466 365614
rect 508702 365378 544466 365614
rect 544702 365378 580466 365614
rect 580702 365378 587342 365614
rect 587578 365378 588670 365614
rect -4746 365366 588670 365378
rect -3826 365354 -3246 365366
rect 4294 365354 4874 365366
rect 40294 365354 40874 365366
rect 76294 365354 76874 365366
rect 112294 365354 112874 365366
rect 148294 365354 148874 365366
rect 184294 365354 184874 365366
rect 220294 365354 220874 365366
rect 256294 365354 256874 365366
rect 292294 365354 292874 365366
rect 328294 365354 328874 365366
rect 364294 365354 364874 365366
rect 400294 365354 400874 365366
rect 436294 365354 436874 365366
rect 472294 365354 472874 365366
rect 508294 365354 508874 365366
rect 544294 365354 544874 365366
rect 580294 365354 580874 365366
rect 587170 365354 587750 365366
rect 238948 363578 248836 363620
rect 238948 363342 238990 363578
rect 239226 363342 248558 363578
rect 248794 363342 248836 363578
rect 238948 363300 248836 363342
rect 268756 363578 345068 363620
rect 268756 363342 268798 363578
rect 269034 363342 344790 363578
rect 345026 363342 345068 363578
rect 268756 363300 345068 363342
rect -1986 362466 -1406 362478
rect 814 362466 1394 362478
rect 36814 362466 37394 362478
rect 72814 362466 73394 362478
rect 108814 362466 109394 362478
rect 144814 362466 145394 362478
rect 180814 362466 181394 362478
rect 216814 362466 217394 362478
rect 252814 362466 253394 362478
rect 288814 362466 289394 362478
rect 324814 362466 325394 362478
rect 360814 362466 361394 362478
rect 396814 362466 397394 362478
rect 432814 362466 433394 362478
rect 468814 362466 469394 362478
rect 504814 362466 505394 362478
rect 540814 362466 541394 362478
rect 576814 362466 577394 362478
rect 585330 362466 585910 362478
rect -2906 362454 586830 362466
rect -2906 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586830 362454
rect -2906 362134 586830 362218
rect -2906 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586830 362134
rect -2906 361886 586830 361898
rect -1986 361874 -1406 361886
rect 814 361874 1394 361886
rect 36814 361874 37394 361886
rect 72814 361874 73394 361886
rect 108814 361874 109394 361886
rect 144814 361874 145394 361886
rect 180814 361874 181394 361886
rect 216814 361874 217394 361886
rect 252814 361874 253394 361886
rect 288814 361874 289394 361886
rect 324814 361874 325394 361886
rect 360814 361874 361394 361886
rect 396814 361874 397394 361886
rect 432814 361874 433394 361886
rect 468814 361874 469394 361886
rect 504814 361874 505394 361886
rect 540814 361874 541394 361886
rect 576814 361874 577394 361886
rect 585330 361874 585910 361886
rect 230668 360858 239268 360900
rect 230668 360622 230710 360858
rect 230946 360622 238990 360858
rect 239226 360622 239268 360858
rect 230668 360580 239268 360622
rect 248516 360858 269076 360900
rect 248516 360622 248558 360858
rect 248794 360622 268798 360858
rect 269034 360622 269076 360858
rect 248516 360580 269076 360622
rect 344748 360858 359788 360900
rect 344748 360622 344790 360858
rect 345026 360622 359510 360858
rect 359746 360622 359788 360858
rect 344748 360580 359788 360622
rect -8426 354906 -7846 354918
rect 29254 354906 29834 354918
rect 65254 354906 65834 354918
rect 101254 354906 101834 354918
rect 137254 354906 137834 354918
rect 173254 354906 173834 354918
rect 209254 354906 209834 354918
rect 245254 354906 245834 354918
rect 281254 354906 281834 354918
rect 317254 354906 317834 354918
rect 353254 354906 353834 354918
rect 389254 354906 389834 354918
rect 425254 354906 425834 354918
rect 461254 354906 461834 354918
rect 497254 354906 497834 354918
rect 533254 354906 533834 354918
rect 569254 354906 569834 354918
rect 591770 354906 592350 354918
rect -8426 354894 592350 354906
rect -8426 354658 -8254 354894
rect -8018 354658 29426 354894
rect 29662 354658 65426 354894
rect 65662 354658 101426 354894
rect 101662 354658 137426 354894
rect 137662 354658 173426 354894
rect 173662 354658 209426 354894
rect 209662 354658 245426 354894
rect 245662 354658 281426 354894
rect 281662 354658 317426 354894
rect 317662 354658 353426 354894
rect 353662 354658 389426 354894
rect 389662 354658 425426 354894
rect 425662 354658 461426 354894
rect 461662 354658 497426 354894
rect 497662 354658 533426 354894
rect 533662 354658 569426 354894
rect 569662 354658 591942 354894
rect 592178 354658 592350 354894
rect -8426 354574 592350 354658
rect -8426 354338 -8254 354574
rect -8018 354338 29426 354574
rect 29662 354338 65426 354574
rect 65662 354338 101426 354574
rect 101662 354338 137426 354574
rect 137662 354338 173426 354574
rect 173662 354338 209426 354574
rect 209662 354338 245426 354574
rect 245662 354338 281426 354574
rect 281662 354338 317426 354574
rect 317662 354338 353426 354574
rect 353662 354338 389426 354574
rect 389662 354338 425426 354574
rect 425662 354338 461426 354574
rect 461662 354338 497426 354574
rect 497662 354338 533426 354574
rect 533662 354338 569426 354574
rect 569662 354338 591942 354574
rect 592178 354338 592350 354574
rect -8426 354326 592350 354338
rect -8426 354314 -7846 354326
rect 29254 354314 29834 354326
rect 65254 354314 65834 354326
rect 101254 354314 101834 354326
rect 137254 354314 137834 354326
rect 173254 354314 173834 354326
rect 209254 354314 209834 354326
rect 245254 354314 245834 354326
rect 281254 354314 281834 354326
rect 317254 354314 317834 354326
rect 353254 354314 353834 354326
rect 389254 354314 389834 354326
rect 425254 354314 425834 354326
rect 461254 354314 461834 354326
rect 497254 354314 497834 354326
rect 533254 354314 533834 354326
rect 569254 354314 569834 354326
rect 591770 354314 592350 354326
rect -6586 351426 -6006 351438
rect 25774 351426 26354 351438
rect 61774 351426 62354 351438
rect 97774 351426 98354 351438
rect 133774 351426 134354 351438
rect 169774 351426 170354 351438
rect 205774 351426 206354 351438
rect 241774 351426 242354 351438
rect 277774 351426 278354 351438
rect 313774 351426 314354 351438
rect 349774 351426 350354 351438
rect 385774 351426 386354 351438
rect 421774 351426 422354 351438
rect 457774 351426 458354 351438
rect 493774 351426 494354 351438
rect 529774 351426 530354 351438
rect 565774 351426 566354 351438
rect 589930 351426 590510 351438
rect -6586 351414 590510 351426
rect -6586 351178 -6414 351414
rect -6178 351178 25946 351414
rect 26182 351178 61946 351414
rect 62182 351178 97946 351414
rect 98182 351178 133946 351414
rect 134182 351178 169946 351414
rect 170182 351178 205946 351414
rect 206182 351178 241946 351414
rect 242182 351178 277946 351414
rect 278182 351178 313946 351414
rect 314182 351178 349946 351414
rect 350182 351178 385946 351414
rect 386182 351178 421946 351414
rect 422182 351178 457946 351414
rect 458182 351178 493946 351414
rect 494182 351178 529946 351414
rect 530182 351178 565946 351414
rect 566182 351178 590102 351414
rect 590338 351178 590510 351414
rect -6586 351094 590510 351178
rect -6586 350858 -6414 351094
rect -6178 350858 25946 351094
rect 26182 350858 61946 351094
rect 62182 350858 97946 351094
rect 98182 350858 133946 351094
rect 134182 350858 169946 351094
rect 170182 350858 205946 351094
rect 206182 350858 241946 351094
rect 242182 350858 277946 351094
rect 278182 350858 313946 351094
rect 314182 350858 349946 351094
rect 350182 350858 385946 351094
rect 386182 350858 421946 351094
rect 422182 350858 457946 351094
rect 458182 350858 493946 351094
rect 494182 350858 529946 351094
rect 530182 350858 565946 351094
rect 566182 350858 590102 351094
rect 590338 350858 590510 351094
rect -6586 350846 590510 350858
rect -6586 350834 -6006 350846
rect 25774 350834 26354 350846
rect 61774 350834 62354 350846
rect 97774 350834 98354 350846
rect 133774 350834 134354 350846
rect 169774 350834 170354 350846
rect 205774 350834 206354 350846
rect 241774 350834 242354 350846
rect 277774 350834 278354 350846
rect 313774 350834 314354 350846
rect 349774 350834 350354 350846
rect 385774 350834 386354 350846
rect 421774 350834 422354 350846
rect 457774 350834 458354 350846
rect 493774 350834 494354 350846
rect 529774 350834 530354 350846
rect 565774 350834 566354 350846
rect 589930 350834 590510 350846
rect -4746 347946 -4166 347958
rect 22294 347946 22874 347958
rect 58294 347946 58874 347958
rect 94294 347946 94874 347958
rect 130294 347946 130874 347958
rect 166294 347946 166874 347958
rect 202294 347946 202874 347958
rect 238294 347946 238874 347958
rect 274294 347946 274874 347958
rect 310294 347946 310874 347958
rect 346294 347946 346874 347958
rect 382294 347946 382874 347958
rect 418294 347946 418874 347958
rect 454294 347946 454874 347958
rect 490294 347946 490874 347958
rect 526294 347946 526874 347958
rect 562294 347946 562874 347958
rect 588090 347946 588670 347958
rect -4746 347934 588670 347946
rect -4746 347698 -4574 347934
rect -4338 347698 22466 347934
rect 22702 347698 58466 347934
rect 58702 347698 94466 347934
rect 94702 347698 130466 347934
rect 130702 347698 166466 347934
rect 166702 347698 202466 347934
rect 202702 347698 238466 347934
rect 238702 347698 274466 347934
rect 274702 347698 310466 347934
rect 310702 347698 346466 347934
rect 346702 347698 382466 347934
rect 382702 347698 418466 347934
rect 418702 347698 454466 347934
rect 454702 347698 490466 347934
rect 490702 347698 526466 347934
rect 526702 347698 562466 347934
rect 562702 347698 588262 347934
rect 588498 347698 588670 347934
rect -4746 347614 588670 347698
rect -4746 347378 -4574 347614
rect -4338 347378 22466 347614
rect 22702 347378 58466 347614
rect 58702 347378 94466 347614
rect 94702 347378 130466 347614
rect 130702 347378 166466 347614
rect 166702 347378 202466 347614
rect 202702 347378 238466 347614
rect 238702 347378 274466 347614
rect 274702 347378 310466 347614
rect 310702 347378 346466 347614
rect 346702 347378 382466 347614
rect 382702 347378 418466 347614
rect 418702 347378 454466 347614
rect 454702 347378 490466 347614
rect 490702 347378 526466 347614
rect 526702 347378 562466 347614
rect 562702 347378 588262 347614
rect 588498 347378 588670 347614
rect -4746 347366 588670 347378
rect -4746 347354 -4166 347366
rect 22294 347354 22874 347366
rect 58294 347354 58874 347366
rect 94294 347354 94874 347366
rect 130294 347354 130874 347366
rect 166294 347354 166874 347366
rect 202294 347354 202874 347366
rect 238294 347354 238874 347366
rect 274294 347354 274874 347366
rect 310294 347354 310874 347366
rect 346294 347354 346874 347366
rect 382294 347354 382874 347366
rect 418294 347354 418874 347366
rect 454294 347354 454874 347366
rect 490294 347354 490874 347366
rect 526294 347354 526874 347366
rect 562294 347354 562874 347366
rect 588090 347354 588670 347366
rect -2906 344466 -2326 344478
rect 18814 344466 19394 344478
rect 54814 344466 55394 344478
rect 90814 344466 91394 344478
rect 126814 344466 127394 344478
rect 162814 344466 163394 344478
rect 198814 344466 199394 344478
rect 234814 344466 235394 344478
rect 270814 344466 271394 344478
rect 306814 344466 307394 344478
rect 342814 344466 343394 344478
rect 378814 344466 379394 344478
rect 414814 344466 415394 344478
rect 450814 344466 451394 344478
rect 486814 344466 487394 344478
rect 522814 344466 523394 344478
rect 558814 344466 559394 344478
rect 586250 344466 586830 344478
rect -2906 344454 586830 344466
rect -2906 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586830 344454
rect -2906 344134 586830 344218
rect -2906 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586830 344134
rect -2906 343886 586830 343898
rect -2906 343874 -2326 343886
rect 18814 343874 19394 343886
rect 54814 343874 55394 343886
rect 90814 343874 91394 343886
rect 126814 343874 127394 343886
rect 162814 343874 163394 343886
rect 198814 343874 199394 343886
rect 234814 343874 235394 343886
rect 270814 343874 271394 343886
rect 306814 343874 307394 343886
rect 342814 343874 343394 343886
rect 378814 343874 379394 343886
rect 414814 343874 415394 343886
rect 450814 343874 451394 343886
rect 486814 343874 487394 343886
rect 522814 343874 523394 343886
rect 558814 343874 559394 343886
rect 586250 343874 586830 343886
rect -7506 336906 -6926 336918
rect 11254 336906 11834 336918
rect 47254 336906 47834 336918
rect 83254 336906 83834 336918
rect 119254 336906 119834 336918
rect 155254 336906 155834 336918
rect 191254 336906 191834 336918
rect 227254 336906 227834 336918
rect 263254 336906 263834 336918
rect 299254 336906 299834 336918
rect 335254 336906 335834 336918
rect 371254 336906 371834 336918
rect 407254 336906 407834 336918
rect 443254 336906 443834 336918
rect 479254 336906 479834 336918
rect 515254 336906 515834 336918
rect 551254 336906 551834 336918
rect 590850 336906 591430 336918
rect -8426 336894 592350 336906
rect -8426 336658 -7334 336894
rect -7098 336658 11426 336894
rect 11662 336658 47426 336894
rect 47662 336658 83426 336894
rect 83662 336658 119426 336894
rect 119662 336658 155426 336894
rect 155662 336658 191426 336894
rect 191662 336658 227426 336894
rect 227662 336658 263426 336894
rect 263662 336658 299426 336894
rect 299662 336658 335426 336894
rect 335662 336658 371426 336894
rect 371662 336658 407426 336894
rect 407662 336658 443426 336894
rect 443662 336658 479426 336894
rect 479662 336658 515426 336894
rect 515662 336658 551426 336894
rect 551662 336658 591022 336894
rect 591258 336658 592350 336894
rect -8426 336574 592350 336658
rect -8426 336338 -7334 336574
rect -7098 336338 11426 336574
rect 11662 336338 47426 336574
rect 47662 336338 83426 336574
rect 83662 336338 119426 336574
rect 119662 336338 155426 336574
rect 155662 336338 191426 336574
rect 191662 336338 227426 336574
rect 227662 336338 263426 336574
rect 263662 336338 299426 336574
rect 299662 336338 335426 336574
rect 335662 336338 371426 336574
rect 371662 336338 407426 336574
rect 407662 336338 443426 336574
rect 443662 336338 479426 336574
rect 479662 336338 515426 336574
rect 515662 336338 551426 336574
rect 551662 336338 591022 336574
rect 591258 336338 592350 336574
rect -8426 336326 592350 336338
rect -7506 336314 -6926 336326
rect 11254 336314 11834 336326
rect 47254 336314 47834 336326
rect 83254 336314 83834 336326
rect 119254 336314 119834 336326
rect 155254 336314 155834 336326
rect 191254 336314 191834 336326
rect 227254 336314 227834 336326
rect 263254 336314 263834 336326
rect 299254 336314 299834 336326
rect 335254 336314 335834 336326
rect 371254 336314 371834 336326
rect 407254 336314 407834 336326
rect 443254 336314 443834 336326
rect 479254 336314 479834 336326
rect 515254 336314 515834 336326
rect 551254 336314 551834 336326
rect 590850 336314 591430 336326
rect -5666 333426 -5086 333438
rect 7774 333426 8354 333438
rect 43774 333426 44354 333438
rect 79774 333426 80354 333438
rect 115774 333426 116354 333438
rect 151774 333426 152354 333438
rect 187774 333426 188354 333438
rect 223774 333426 224354 333438
rect 259774 333426 260354 333438
rect 295774 333426 296354 333438
rect 331774 333426 332354 333438
rect 367774 333426 368354 333438
rect 403774 333426 404354 333438
rect 439774 333426 440354 333438
rect 475774 333426 476354 333438
rect 511774 333426 512354 333438
rect 547774 333426 548354 333438
rect 589010 333426 589590 333438
rect -6586 333414 590510 333426
rect -6586 333178 -5494 333414
rect -5258 333178 7946 333414
rect 8182 333178 43946 333414
rect 44182 333178 79946 333414
rect 80182 333178 115946 333414
rect 116182 333178 151946 333414
rect 152182 333178 187946 333414
rect 188182 333178 223946 333414
rect 224182 333178 259946 333414
rect 260182 333178 295946 333414
rect 296182 333178 331946 333414
rect 332182 333178 367946 333414
rect 368182 333178 403946 333414
rect 404182 333178 439946 333414
rect 440182 333178 475946 333414
rect 476182 333178 511946 333414
rect 512182 333178 547946 333414
rect 548182 333178 589182 333414
rect 589418 333178 590510 333414
rect -6586 333094 590510 333178
rect -6586 332858 -5494 333094
rect -5258 332858 7946 333094
rect 8182 332858 43946 333094
rect 44182 332858 79946 333094
rect 80182 332858 115946 333094
rect 116182 332858 151946 333094
rect 152182 332858 187946 333094
rect 188182 332858 223946 333094
rect 224182 332858 259946 333094
rect 260182 332858 295946 333094
rect 296182 332858 331946 333094
rect 332182 332858 367946 333094
rect 368182 332858 403946 333094
rect 404182 332858 439946 333094
rect 440182 332858 475946 333094
rect 476182 332858 511946 333094
rect 512182 332858 547946 333094
rect 548182 332858 589182 333094
rect 589418 332858 590510 333094
rect -6586 332846 590510 332858
rect -5666 332834 -5086 332846
rect 7774 332834 8354 332846
rect 43774 332834 44354 332846
rect 79774 332834 80354 332846
rect 115774 332834 116354 332846
rect 151774 332834 152354 332846
rect 187774 332834 188354 332846
rect 223774 332834 224354 332846
rect 259774 332834 260354 332846
rect 295774 332834 296354 332846
rect 331774 332834 332354 332846
rect 367774 332834 368354 332846
rect 403774 332834 404354 332846
rect 439774 332834 440354 332846
rect 475774 332834 476354 332846
rect 511774 332834 512354 332846
rect 547774 332834 548354 332846
rect 589010 332834 589590 332846
rect -3826 329946 -3246 329958
rect 4294 329946 4874 329958
rect 40294 329946 40874 329958
rect 76294 329946 76874 329958
rect 112294 329946 112874 329958
rect 148294 329946 148874 329958
rect 184294 329946 184874 329958
rect 220294 329946 220874 329958
rect 256294 329946 256874 329958
rect 292294 329946 292874 329958
rect 328294 329946 328874 329958
rect 364294 329946 364874 329958
rect 400294 329946 400874 329958
rect 436294 329946 436874 329958
rect 472294 329946 472874 329958
rect 508294 329946 508874 329958
rect 544294 329946 544874 329958
rect 580294 329946 580874 329958
rect 587170 329946 587750 329958
rect -4746 329934 588670 329946
rect -4746 329698 -3654 329934
rect -3418 329698 4466 329934
rect 4702 329698 40466 329934
rect 40702 329698 76466 329934
rect 76702 329698 112466 329934
rect 112702 329698 148466 329934
rect 148702 329698 184466 329934
rect 184702 329698 220466 329934
rect 220702 329698 256466 329934
rect 256702 329698 292466 329934
rect 292702 329698 328466 329934
rect 328702 329698 364466 329934
rect 364702 329698 400466 329934
rect 400702 329698 436466 329934
rect 436702 329698 472466 329934
rect 472702 329698 508466 329934
rect 508702 329698 544466 329934
rect 544702 329698 580466 329934
rect 580702 329698 587342 329934
rect 587578 329698 588670 329934
rect -4746 329614 588670 329698
rect -4746 329378 -3654 329614
rect -3418 329378 4466 329614
rect 4702 329378 40466 329614
rect 40702 329378 76466 329614
rect 76702 329378 112466 329614
rect 112702 329378 148466 329614
rect 148702 329378 184466 329614
rect 184702 329378 220466 329614
rect 220702 329378 256466 329614
rect 256702 329378 292466 329614
rect 292702 329378 328466 329614
rect 328702 329378 364466 329614
rect 364702 329378 400466 329614
rect 400702 329378 436466 329614
rect 436702 329378 472466 329614
rect 472702 329378 508466 329614
rect 508702 329378 544466 329614
rect 544702 329378 580466 329614
rect 580702 329378 587342 329614
rect 587578 329378 588670 329614
rect -4746 329366 588670 329378
rect -3826 329354 -3246 329366
rect 4294 329354 4874 329366
rect 40294 329354 40874 329366
rect 76294 329354 76874 329366
rect 112294 329354 112874 329366
rect 148294 329354 148874 329366
rect 184294 329354 184874 329366
rect 220294 329354 220874 329366
rect 256294 329354 256874 329366
rect 292294 329354 292874 329366
rect 328294 329354 328874 329366
rect 364294 329354 364874 329366
rect 400294 329354 400874 329366
rect 436294 329354 436874 329366
rect 472294 329354 472874 329366
rect 508294 329354 508874 329366
rect 544294 329354 544874 329366
rect 580294 329354 580874 329366
rect 587170 329354 587750 329366
rect -1986 326466 -1406 326478
rect 814 326466 1394 326478
rect 36814 326466 37394 326478
rect 72814 326466 73394 326478
rect 108814 326466 109394 326478
rect 144814 326466 145394 326478
rect 180814 326466 181394 326478
rect 216814 326466 217394 326478
rect 252814 326466 253394 326478
rect 288814 326466 289394 326478
rect 324814 326466 325394 326478
rect 360814 326466 361394 326478
rect 396814 326466 397394 326478
rect 432814 326466 433394 326478
rect 468814 326466 469394 326478
rect 504814 326466 505394 326478
rect 540814 326466 541394 326478
rect 576814 326466 577394 326478
rect 585330 326466 585910 326478
rect -2906 326454 586830 326466
rect -2906 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586830 326454
rect -2906 326134 586830 326218
rect -2906 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586830 326134
rect -2906 325886 586830 325898
rect -1986 325874 -1406 325886
rect 814 325874 1394 325886
rect 36814 325874 37394 325886
rect 72814 325874 73394 325886
rect 108814 325874 109394 325886
rect 144814 325874 145394 325886
rect 180814 325874 181394 325886
rect 216814 325874 217394 325886
rect 252814 325874 253394 325886
rect 288814 325874 289394 325886
rect 324814 325874 325394 325886
rect 360814 325874 361394 325886
rect 396814 325874 397394 325886
rect 432814 325874 433394 325886
rect 468814 325874 469394 325886
rect 504814 325874 505394 325886
rect 540814 325874 541394 325886
rect 576814 325874 577394 325886
rect 585330 325874 585910 325886
rect -8426 318906 -7846 318918
rect 29254 318906 29834 318918
rect 65254 318906 65834 318918
rect 101254 318906 101834 318918
rect 137254 318906 137834 318918
rect 173254 318906 173834 318918
rect 209254 318906 209834 318918
rect 245254 318906 245834 318918
rect 281254 318906 281834 318918
rect 317254 318906 317834 318918
rect 353254 318906 353834 318918
rect 389254 318906 389834 318918
rect 425254 318906 425834 318918
rect 461254 318906 461834 318918
rect 497254 318906 497834 318918
rect 533254 318906 533834 318918
rect 569254 318906 569834 318918
rect 591770 318906 592350 318918
rect -8426 318894 592350 318906
rect -8426 318658 -8254 318894
rect -8018 318658 29426 318894
rect 29662 318658 65426 318894
rect 65662 318658 101426 318894
rect 101662 318658 137426 318894
rect 137662 318658 173426 318894
rect 173662 318658 209426 318894
rect 209662 318658 245426 318894
rect 245662 318658 281426 318894
rect 281662 318658 317426 318894
rect 317662 318658 353426 318894
rect 353662 318658 389426 318894
rect 389662 318658 425426 318894
rect 425662 318658 461426 318894
rect 461662 318658 497426 318894
rect 497662 318658 533426 318894
rect 533662 318658 569426 318894
rect 569662 318658 591942 318894
rect 592178 318658 592350 318894
rect -8426 318574 592350 318658
rect -8426 318338 -8254 318574
rect -8018 318338 29426 318574
rect 29662 318338 65426 318574
rect 65662 318338 101426 318574
rect 101662 318338 137426 318574
rect 137662 318338 173426 318574
rect 173662 318338 209426 318574
rect 209662 318338 245426 318574
rect 245662 318338 281426 318574
rect 281662 318338 317426 318574
rect 317662 318338 353426 318574
rect 353662 318338 389426 318574
rect 389662 318338 425426 318574
rect 425662 318338 461426 318574
rect 461662 318338 497426 318574
rect 497662 318338 533426 318574
rect 533662 318338 569426 318574
rect 569662 318338 591942 318574
rect 592178 318338 592350 318574
rect -8426 318326 592350 318338
rect -8426 318314 -7846 318326
rect 29254 318314 29834 318326
rect 65254 318314 65834 318326
rect 101254 318314 101834 318326
rect 137254 318314 137834 318326
rect 173254 318314 173834 318326
rect 209254 318314 209834 318326
rect 245254 318314 245834 318326
rect 281254 318314 281834 318326
rect 317254 318314 317834 318326
rect 353254 318314 353834 318326
rect 389254 318314 389834 318326
rect 425254 318314 425834 318326
rect 461254 318314 461834 318326
rect 497254 318314 497834 318326
rect 533254 318314 533834 318326
rect 569254 318314 569834 318326
rect 591770 318314 592350 318326
rect -6586 315426 -6006 315438
rect 25774 315426 26354 315438
rect 61774 315426 62354 315438
rect 97774 315426 98354 315438
rect 133774 315426 134354 315438
rect 169774 315426 170354 315438
rect 205774 315426 206354 315438
rect 241774 315426 242354 315438
rect 277774 315426 278354 315438
rect 313774 315426 314354 315438
rect 349774 315426 350354 315438
rect 385774 315426 386354 315438
rect 421774 315426 422354 315438
rect 457774 315426 458354 315438
rect 493774 315426 494354 315438
rect 529774 315426 530354 315438
rect 565774 315426 566354 315438
rect 589930 315426 590510 315438
rect -6586 315414 590510 315426
rect -6586 315178 -6414 315414
rect -6178 315178 25946 315414
rect 26182 315178 61946 315414
rect 62182 315178 97946 315414
rect 98182 315178 133946 315414
rect 134182 315178 169946 315414
rect 170182 315178 205946 315414
rect 206182 315178 241946 315414
rect 242182 315178 277946 315414
rect 278182 315178 313946 315414
rect 314182 315178 349946 315414
rect 350182 315178 385946 315414
rect 386182 315178 421946 315414
rect 422182 315178 457946 315414
rect 458182 315178 493946 315414
rect 494182 315178 529946 315414
rect 530182 315178 565946 315414
rect 566182 315178 590102 315414
rect 590338 315178 590510 315414
rect -6586 315094 590510 315178
rect -6586 314858 -6414 315094
rect -6178 314858 25946 315094
rect 26182 314858 61946 315094
rect 62182 314858 97946 315094
rect 98182 314858 133946 315094
rect 134182 314858 169946 315094
rect 170182 314858 205946 315094
rect 206182 314858 241946 315094
rect 242182 314858 277946 315094
rect 278182 314858 313946 315094
rect 314182 314858 349946 315094
rect 350182 314858 385946 315094
rect 386182 314858 421946 315094
rect 422182 314858 457946 315094
rect 458182 314858 493946 315094
rect 494182 314858 529946 315094
rect 530182 314858 565946 315094
rect 566182 314858 590102 315094
rect 590338 314858 590510 315094
rect -6586 314846 590510 314858
rect -6586 314834 -6006 314846
rect 25774 314834 26354 314846
rect 61774 314834 62354 314846
rect 97774 314834 98354 314846
rect 133774 314834 134354 314846
rect 169774 314834 170354 314846
rect 205774 314834 206354 314846
rect 241774 314834 242354 314846
rect 277774 314834 278354 314846
rect 313774 314834 314354 314846
rect 349774 314834 350354 314846
rect 385774 314834 386354 314846
rect 421774 314834 422354 314846
rect 457774 314834 458354 314846
rect 493774 314834 494354 314846
rect 529774 314834 530354 314846
rect 565774 314834 566354 314846
rect 589930 314834 590510 314846
rect -4746 311946 -4166 311958
rect 22294 311946 22874 311958
rect 58294 311946 58874 311958
rect 94294 311946 94874 311958
rect 130294 311946 130874 311958
rect 166294 311946 166874 311958
rect 202294 311946 202874 311958
rect 238294 311946 238874 311958
rect 274294 311946 274874 311958
rect 310294 311946 310874 311958
rect 346294 311946 346874 311958
rect 382294 311946 382874 311958
rect 418294 311946 418874 311958
rect 454294 311946 454874 311958
rect 490294 311946 490874 311958
rect 526294 311946 526874 311958
rect 562294 311946 562874 311958
rect 588090 311946 588670 311958
rect -4746 311934 588670 311946
rect -4746 311698 -4574 311934
rect -4338 311698 22466 311934
rect 22702 311698 58466 311934
rect 58702 311698 94466 311934
rect 94702 311698 130466 311934
rect 130702 311698 166466 311934
rect 166702 311698 202466 311934
rect 202702 311698 238466 311934
rect 238702 311698 274466 311934
rect 274702 311698 310466 311934
rect 310702 311698 346466 311934
rect 346702 311698 382466 311934
rect 382702 311698 418466 311934
rect 418702 311698 454466 311934
rect 454702 311698 490466 311934
rect 490702 311698 526466 311934
rect 526702 311698 562466 311934
rect 562702 311698 588262 311934
rect 588498 311698 588670 311934
rect -4746 311614 588670 311698
rect -4746 311378 -4574 311614
rect -4338 311378 22466 311614
rect 22702 311378 58466 311614
rect 58702 311378 94466 311614
rect 94702 311378 130466 311614
rect 130702 311378 166466 311614
rect 166702 311378 202466 311614
rect 202702 311378 238466 311614
rect 238702 311378 274466 311614
rect 274702 311378 310466 311614
rect 310702 311378 346466 311614
rect 346702 311378 382466 311614
rect 382702 311378 418466 311614
rect 418702 311378 454466 311614
rect 454702 311378 490466 311614
rect 490702 311378 526466 311614
rect 526702 311378 562466 311614
rect 562702 311378 588262 311614
rect 588498 311378 588670 311614
rect -4746 311366 588670 311378
rect -4746 311354 -4166 311366
rect 22294 311354 22874 311366
rect 58294 311354 58874 311366
rect 94294 311354 94874 311366
rect 130294 311354 130874 311366
rect 166294 311354 166874 311366
rect 202294 311354 202874 311366
rect 238294 311354 238874 311366
rect 274294 311354 274874 311366
rect 310294 311354 310874 311366
rect 346294 311354 346874 311366
rect 382294 311354 382874 311366
rect 418294 311354 418874 311366
rect 454294 311354 454874 311366
rect 490294 311354 490874 311366
rect 526294 311354 526874 311366
rect 562294 311354 562874 311366
rect 588090 311354 588670 311366
rect -2906 308466 -2326 308478
rect 18814 308466 19394 308478
rect 54814 308466 55394 308478
rect 90814 308466 91394 308478
rect 126814 308466 127394 308478
rect 162814 308466 163394 308478
rect 198814 308466 199394 308478
rect 234814 308466 235394 308478
rect 270814 308466 271394 308478
rect 306814 308466 307394 308478
rect 342814 308466 343394 308478
rect 378814 308466 379394 308478
rect 414814 308466 415394 308478
rect 450814 308466 451394 308478
rect 486814 308466 487394 308478
rect 522814 308466 523394 308478
rect 558814 308466 559394 308478
rect 586250 308466 586830 308478
rect -2906 308454 586830 308466
rect -2906 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586830 308454
rect -2906 308134 586830 308218
rect -2906 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586830 308134
rect -2906 307886 586830 307898
rect -2906 307874 -2326 307886
rect 18814 307874 19394 307886
rect 54814 307874 55394 307886
rect 90814 307874 91394 307886
rect 126814 307874 127394 307886
rect 162814 307874 163394 307886
rect 198814 307874 199394 307886
rect 234814 307874 235394 307886
rect 270814 307874 271394 307886
rect 306814 307874 307394 307886
rect 342814 307874 343394 307886
rect 378814 307874 379394 307886
rect 414814 307874 415394 307886
rect 450814 307874 451394 307886
rect 486814 307874 487394 307886
rect 522814 307874 523394 307886
rect 558814 307874 559394 307886
rect 586250 307874 586830 307886
rect -7506 300906 -6926 300918
rect 11254 300906 11834 300918
rect 47254 300906 47834 300918
rect 83254 300906 83834 300918
rect 119254 300906 119834 300918
rect 155254 300906 155834 300918
rect 191254 300906 191834 300918
rect 227254 300906 227834 300918
rect 263254 300906 263834 300918
rect 299254 300906 299834 300918
rect 335254 300906 335834 300918
rect 371254 300906 371834 300918
rect 407254 300906 407834 300918
rect 443254 300906 443834 300918
rect 479254 300906 479834 300918
rect 515254 300906 515834 300918
rect 551254 300906 551834 300918
rect 590850 300906 591430 300918
rect -8426 300894 592350 300906
rect -8426 300658 -7334 300894
rect -7098 300658 11426 300894
rect 11662 300658 47426 300894
rect 47662 300658 83426 300894
rect 83662 300658 119426 300894
rect 119662 300658 155426 300894
rect 155662 300658 191426 300894
rect 191662 300658 227426 300894
rect 227662 300658 263426 300894
rect 263662 300658 299426 300894
rect 299662 300658 335426 300894
rect 335662 300658 371426 300894
rect 371662 300658 407426 300894
rect 407662 300658 443426 300894
rect 443662 300658 479426 300894
rect 479662 300658 515426 300894
rect 515662 300658 551426 300894
rect 551662 300658 591022 300894
rect 591258 300658 592350 300894
rect -8426 300574 592350 300658
rect -8426 300338 -7334 300574
rect -7098 300338 11426 300574
rect 11662 300338 47426 300574
rect 47662 300338 83426 300574
rect 83662 300338 119426 300574
rect 119662 300338 155426 300574
rect 155662 300338 191426 300574
rect 191662 300338 227426 300574
rect 227662 300338 263426 300574
rect 263662 300338 299426 300574
rect 299662 300338 335426 300574
rect 335662 300338 371426 300574
rect 371662 300338 407426 300574
rect 407662 300338 443426 300574
rect 443662 300338 479426 300574
rect 479662 300338 515426 300574
rect 515662 300338 551426 300574
rect 551662 300338 591022 300574
rect 591258 300338 592350 300574
rect -8426 300326 592350 300338
rect -7506 300314 -6926 300326
rect 11254 300314 11834 300326
rect 47254 300314 47834 300326
rect 83254 300314 83834 300326
rect 119254 300314 119834 300326
rect 155254 300314 155834 300326
rect 191254 300314 191834 300326
rect 227254 300314 227834 300326
rect 263254 300314 263834 300326
rect 299254 300314 299834 300326
rect 335254 300314 335834 300326
rect 371254 300314 371834 300326
rect 407254 300314 407834 300326
rect 443254 300314 443834 300326
rect 479254 300314 479834 300326
rect 515254 300314 515834 300326
rect 551254 300314 551834 300326
rect 590850 300314 591430 300326
rect -5666 297426 -5086 297438
rect 7774 297426 8354 297438
rect 43774 297426 44354 297438
rect 79774 297426 80354 297438
rect 115774 297426 116354 297438
rect 151774 297426 152354 297438
rect 187774 297426 188354 297438
rect 223774 297426 224354 297438
rect 259774 297426 260354 297438
rect 295774 297426 296354 297438
rect 331774 297426 332354 297438
rect 367774 297426 368354 297438
rect 403774 297426 404354 297438
rect 439774 297426 440354 297438
rect 475774 297426 476354 297438
rect 511774 297426 512354 297438
rect 547774 297426 548354 297438
rect 589010 297426 589590 297438
rect -6586 297414 590510 297426
rect -6586 297178 -5494 297414
rect -5258 297178 7946 297414
rect 8182 297178 43946 297414
rect 44182 297178 79946 297414
rect 80182 297178 115946 297414
rect 116182 297178 151946 297414
rect 152182 297178 187946 297414
rect 188182 297178 223946 297414
rect 224182 297178 259946 297414
rect 260182 297178 295946 297414
rect 296182 297178 331946 297414
rect 332182 297178 367946 297414
rect 368182 297178 403946 297414
rect 404182 297178 439946 297414
rect 440182 297178 475946 297414
rect 476182 297178 511946 297414
rect 512182 297178 547946 297414
rect 548182 297178 589182 297414
rect 589418 297178 590510 297414
rect -6586 297094 590510 297178
rect -6586 296858 -5494 297094
rect -5258 296858 7946 297094
rect 8182 296858 43946 297094
rect 44182 296858 79946 297094
rect 80182 296858 115946 297094
rect 116182 296858 151946 297094
rect 152182 296858 187946 297094
rect 188182 296858 223946 297094
rect 224182 296858 259946 297094
rect 260182 296858 295946 297094
rect 296182 296858 331946 297094
rect 332182 296858 367946 297094
rect 368182 296858 403946 297094
rect 404182 296858 439946 297094
rect 440182 296858 475946 297094
rect 476182 296858 511946 297094
rect 512182 296858 547946 297094
rect 548182 296858 589182 297094
rect 589418 296858 590510 297094
rect -6586 296846 590510 296858
rect -5666 296834 -5086 296846
rect 7774 296834 8354 296846
rect 43774 296834 44354 296846
rect 79774 296834 80354 296846
rect 115774 296834 116354 296846
rect 151774 296834 152354 296846
rect 187774 296834 188354 296846
rect 223774 296834 224354 296846
rect 259774 296834 260354 296846
rect 295774 296834 296354 296846
rect 331774 296834 332354 296846
rect 367774 296834 368354 296846
rect 403774 296834 404354 296846
rect 439774 296834 440354 296846
rect 475774 296834 476354 296846
rect 511774 296834 512354 296846
rect 547774 296834 548354 296846
rect 589010 296834 589590 296846
rect -3826 293946 -3246 293958
rect 4294 293946 4874 293958
rect 40294 293946 40874 293958
rect 76294 293946 76874 293958
rect 112294 293946 112874 293958
rect 148294 293946 148874 293958
rect 184294 293946 184874 293958
rect 220294 293946 220874 293958
rect 256294 293946 256874 293958
rect 292294 293946 292874 293958
rect 328294 293946 328874 293958
rect 364294 293946 364874 293958
rect 400294 293946 400874 293958
rect 436294 293946 436874 293958
rect 472294 293946 472874 293958
rect 508294 293946 508874 293958
rect 544294 293946 544874 293958
rect 580294 293946 580874 293958
rect 587170 293946 587750 293958
rect -4746 293934 588670 293946
rect -4746 293698 -3654 293934
rect -3418 293698 4466 293934
rect 4702 293698 40466 293934
rect 40702 293698 76466 293934
rect 76702 293698 112466 293934
rect 112702 293698 148466 293934
rect 148702 293698 184466 293934
rect 184702 293698 220466 293934
rect 220702 293698 256466 293934
rect 256702 293698 292466 293934
rect 292702 293698 328466 293934
rect 328702 293698 364466 293934
rect 364702 293698 400466 293934
rect 400702 293698 436466 293934
rect 436702 293698 472466 293934
rect 472702 293698 508466 293934
rect 508702 293698 544466 293934
rect 544702 293698 580466 293934
rect 580702 293698 587342 293934
rect 587578 293698 588670 293934
rect -4746 293614 588670 293698
rect -4746 293378 -3654 293614
rect -3418 293378 4466 293614
rect 4702 293378 40466 293614
rect 40702 293378 76466 293614
rect 76702 293378 112466 293614
rect 112702 293378 148466 293614
rect 148702 293378 184466 293614
rect 184702 293378 220466 293614
rect 220702 293378 256466 293614
rect 256702 293378 292466 293614
rect 292702 293378 328466 293614
rect 328702 293378 364466 293614
rect 364702 293378 400466 293614
rect 400702 293378 436466 293614
rect 436702 293378 472466 293614
rect 472702 293378 508466 293614
rect 508702 293378 544466 293614
rect 544702 293378 580466 293614
rect 580702 293378 587342 293614
rect 587578 293378 588670 293614
rect -4746 293366 588670 293378
rect -3826 293354 -3246 293366
rect 4294 293354 4874 293366
rect 40294 293354 40874 293366
rect 76294 293354 76874 293366
rect 112294 293354 112874 293366
rect 148294 293354 148874 293366
rect 184294 293354 184874 293366
rect 220294 293354 220874 293366
rect 256294 293354 256874 293366
rect 292294 293354 292874 293366
rect 328294 293354 328874 293366
rect 364294 293354 364874 293366
rect 400294 293354 400874 293366
rect 436294 293354 436874 293366
rect 472294 293354 472874 293366
rect 508294 293354 508874 293366
rect 544294 293354 544874 293366
rect 580294 293354 580874 293366
rect 587170 293354 587750 293366
rect -1986 290466 -1406 290478
rect 814 290466 1394 290478
rect 36814 290466 37394 290478
rect 72814 290466 73394 290478
rect 108814 290466 109394 290478
rect 144814 290466 145394 290478
rect 180814 290466 181394 290478
rect 216814 290466 217394 290478
rect 252814 290466 253394 290478
rect 288814 290466 289394 290478
rect 324814 290466 325394 290478
rect 360814 290466 361394 290478
rect 396814 290466 397394 290478
rect 432814 290466 433394 290478
rect 468814 290466 469394 290478
rect 504814 290466 505394 290478
rect 540814 290466 541394 290478
rect 576814 290466 577394 290478
rect 585330 290466 585910 290478
rect -2906 290454 586830 290466
rect -2906 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586830 290454
rect -2906 290134 586830 290218
rect -2906 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586830 290134
rect -2906 289886 586830 289898
rect -1986 289874 -1406 289886
rect 814 289874 1394 289886
rect 36814 289874 37394 289886
rect 72814 289874 73394 289886
rect 108814 289874 109394 289886
rect 144814 289874 145394 289886
rect 180814 289874 181394 289886
rect 216814 289874 217394 289886
rect 252814 289874 253394 289886
rect 288814 289874 289394 289886
rect 324814 289874 325394 289886
rect 360814 289874 361394 289886
rect 396814 289874 397394 289886
rect 432814 289874 433394 289886
rect 468814 289874 469394 289886
rect 504814 289874 505394 289886
rect 540814 289874 541394 289886
rect 576814 289874 577394 289886
rect 585330 289874 585910 289886
rect -8426 282906 -7846 282918
rect 29254 282906 29834 282918
rect 65254 282906 65834 282918
rect 101254 282906 101834 282918
rect 137254 282906 137834 282918
rect 173254 282906 173834 282918
rect 209254 282906 209834 282918
rect 245254 282906 245834 282918
rect 281254 282906 281834 282918
rect 317254 282906 317834 282918
rect 353254 282906 353834 282918
rect 389254 282906 389834 282918
rect 425254 282906 425834 282918
rect 461254 282906 461834 282918
rect 497254 282906 497834 282918
rect 533254 282906 533834 282918
rect 569254 282906 569834 282918
rect 591770 282906 592350 282918
rect -8426 282894 592350 282906
rect -8426 282658 -8254 282894
rect -8018 282658 29426 282894
rect 29662 282658 65426 282894
rect 65662 282658 101426 282894
rect 101662 282658 137426 282894
rect 137662 282658 173426 282894
rect 173662 282658 209426 282894
rect 209662 282658 245426 282894
rect 245662 282658 281426 282894
rect 281662 282658 317426 282894
rect 317662 282658 353426 282894
rect 353662 282658 389426 282894
rect 389662 282658 425426 282894
rect 425662 282658 461426 282894
rect 461662 282658 497426 282894
rect 497662 282658 533426 282894
rect 533662 282658 569426 282894
rect 569662 282658 591942 282894
rect 592178 282658 592350 282894
rect -8426 282574 592350 282658
rect -8426 282338 -8254 282574
rect -8018 282338 29426 282574
rect 29662 282338 65426 282574
rect 65662 282338 101426 282574
rect 101662 282338 137426 282574
rect 137662 282338 173426 282574
rect 173662 282338 209426 282574
rect 209662 282338 245426 282574
rect 245662 282338 281426 282574
rect 281662 282338 317426 282574
rect 317662 282338 353426 282574
rect 353662 282338 389426 282574
rect 389662 282338 425426 282574
rect 425662 282338 461426 282574
rect 461662 282338 497426 282574
rect 497662 282338 533426 282574
rect 533662 282338 569426 282574
rect 569662 282338 591942 282574
rect 592178 282338 592350 282574
rect -8426 282326 592350 282338
rect -8426 282314 -7846 282326
rect 29254 282314 29834 282326
rect 65254 282314 65834 282326
rect 101254 282314 101834 282326
rect 137254 282314 137834 282326
rect 173254 282314 173834 282326
rect 209254 282314 209834 282326
rect 245254 282314 245834 282326
rect 281254 282314 281834 282326
rect 317254 282314 317834 282326
rect 353254 282314 353834 282326
rect 389254 282314 389834 282326
rect 425254 282314 425834 282326
rect 461254 282314 461834 282326
rect 497254 282314 497834 282326
rect 533254 282314 533834 282326
rect 569254 282314 569834 282326
rect 591770 282314 592350 282326
rect -6586 279426 -6006 279438
rect 25774 279426 26354 279438
rect 61774 279426 62354 279438
rect 97774 279426 98354 279438
rect 133774 279426 134354 279438
rect 169774 279426 170354 279438
rect 205774 279426 206354 279438
rect 241774 279426 242354 279438
rect 277774 279426 278354 279438
rect 313774 279426 314354 279438
rect 349774 279426 350354 279438
rect 385774 279426 386354 279438
rect 421774 279426 422354 279438
rect 457774 279426 458354 279438
rect 493774 279426 494354 279438
rect 529774 279426 530354 279438
rect 565774 279426 566354 279438
rect 589930 279426 590510 279438
rect -6586 279414 590510 279426
rect -6586 279178 -6414 279414
rect -6178 279178 25946 279414
rect 26182 279178 61946 279414
rect 62182 279178 97946 279414
rect 98182 279178 133946 279414
rect 134182 279178 169946 279414
rect 170182 279178 205946 279414
rect 206182 279178 241946 279414
rect 242182 279178 277946 279414
rect 278182 279178 313946 279414
rect 314182 279178 349946 279414
rect 350182 279178 385946 279414
rect 386182 279178 421946 279414
rect 422182 279178 457946 279414
rect 458182 279178 493946 279414
rect 494182 279178 529946 279414
rect 530182 279178 565946 279414
rect 566182 279178 590102 279414
rect 590338 279178 590510 279414
rect -6586 279094 590510 279178
rect -6586 278858 -6414 279094
rect -6178 278858 25946 279094
rect 26182 278858 61946 279094
rect 62182 278858 97946 279094
rect 98182 278858 133946 279094
rect 134182 278858 169946 279094
rect 170182 278858 205946 279094
rect 206182 278858 241946 279094
rect 242182 278858 277946 279094
rect 278182 278858 313946 279094
rect 314182 278858 349946 279094
rect 350182 278858 385946 279094
rect 386182 278858 421946 279094
rect 422182 278858 457946 279094
rect 458182 278858 493946 279094
rect 494182 278858 529946 279094
rect 530182 278858 565946 279094
rect 566182 278858 590102 279094
rect 590338 278858 590510 279094
rect -6586 278846 590510 278858
rect -6586 278834 -6006 278846
rect 25774 278834 26354 278846
rect 61774 278834 62354 278846
rect 97774 278834 98354 278846
rect 133774 278834 134354 278846
rect 169774 278834 170354 278846
rect 205774 278834 206354 278846
rect 241774 278834 242354 278846
rect 277774 278834 278354 278846
rect 313774 278834 314354 278846
rect 349774 278834 350354 278846
rect 385774 278834 386354 278846
rect 421774 278834 422354 278846
rect 457774 278834 458354 278846
rect 493774 278834 494354 278846
rect 529774 278834 530354 278846
rect 565774 278834 566354 278846
rect 589930 278834 590510 278846
rect -4746 275946 -4166 275958
rect 22294 275946 22874 275958
rect 58294 275946 58874 275958
rect 94294 275946 94874 275958
rect 130294 275946 130874 275958
rect 166294 275946 166874 275958
rect 202294 275946 202874 275958
rect 238294 275946 238874 275958
rect 274294 275946 274874 275958
rect 310294 275946 310874 275958
rect 346294 275946 346874 275958
rect 382294 275946 382874 275958
rect 418294 275946 418874 275958
rect 454294 275946 454874 275958
rect 490294 275946 490874 275958
rect 526294 275946 526874 275958
rect 562294 275946 562874 275958
rect 588090 275946 588670 275958
rect -4746 275934 588670 275946
rect -4746 275698 -4574 275934
rect -4338 275698 22466 275934
rect 22702 275698 58466 275934
rect 58702 275698 94466 275934
rect 94702 275698 130466 275934
rect 130702 275698 166466 275934
rect 166702 275698 202466 275934
rect 202702 275698 238466 275934
rect 238702 275698 274466 275934
rect 274702 275698 310466 275934
rect 310702 275698 346466 275934
rect 346702 275698 382466 275934
rect 382702 275698 418466 275934
rect 418702 275698 454466 275934
rect 454702 275698 490466 275934
rect 490702 275698 526466 275934
rect 526702 275698 562466 275934
rect 562702 275698 588262 275934
rect 588498 275698 588670 275934
rect -4746 275614 588670 275698
rect -4746 275378 -4574 275614
rect -4338 275378 22466 275614
rect 22702 275378 58466 275614
rect 58702 275378 94466 275614
rect 94702 275378 130466 275614
rect 130702 275378 166466 275614
rect 166702 275378 202466 275614
rect 202702 275378 238466 275614
rect 238702 275378 274466 275614
rect 274702 275378 310466 275614
rect 310702 275378 346466 275614
rect 346702 275378 382466 275614
rect 382702 275378 418466 275614
rect 418702 275378 454466 275614
rect 454702 275378 490466 275614
rect 490702 275378 526466 275614
rect 526702 275378 562466 275614
rect 562702 275378 588262 275614
rect 588498 275378 588670 275614
rect -4746 275366 588670 275378
rect -4746 275354 -4166 275366
rect 22294 275354 22874 275366
rect 58294 275354 58874 275366
rect 94294 275354 94874 275366
rect 130294 275354 130874 275366
rect 166294 275354 166874 275366
rect 202294 275354 202874 275366
rect 238294 275354 238874 275366
rect 274294 275354 274874 275366
rect 310294 275354 310874 275366
rect 346294 275354 346874 275366
rect 382294 275354 382874 275366
rect 418294 275354 418874 275366
rect 454294 275354 454874 275366
rect 490294 275354 490874 275366
rect 526294 275354 526874 275366
rect 562294 275354 562874 275366
rect 588090 275354 588670 275366
rect -2906 272466 -2326 272478
rect 18814 272466 19394 272478
rect 54814 272466 55394 272478
rect 90814 272466 91394 272478
rect 126814 272466 127394 272478
rect 162814 272466 163394 272478
rect 198814 272466 199394 272478
rect 234814 272466 235394 272478
rect 270814 272466 271394 272478
rect 306814 272466 307394 272478
rect 342814 272466 343394 272478
rect 378814 272466 379394 272478
rect 414814 272466 415394 272478
rect 450814 272466 451394 272478
rect 486814 272466 487394 272478
rect 522814 272466 523394 272478
rect 558814 272466 559394 272478
rect 586250 272466 586830 272478
rect -2906 272454 586830 272466
rect -2906 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586830 272454
rect -2906 272134 586830 272218
rect -2906 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586830 272134
rect -2906 271886 586830 271898
rect -2906 271874 -2326 271886
rect 18814 271874 19394 271886
rect 54814 271874 55394 271886
rect 90814 271874 91394 271886
rect 126814 271874 127394 271886
rect 162814 271874 163394 271886
rect 198814 271874 199394 271886
rect 234814 271874 235394 271886
rect 270814 271874 271394 271886
rect 306814 271874 307394 271886
rect 342814 271874 343394 271886
rect 378814 271874 379394 271886
rect 414814 271874 415394 271886
rect 450814 271874 451394 271886
rect 486814 271874 487394 271886
rect 522814 271874 523394 271886
rect 558814 271874 559394 271886
rect 586250 271874 586830 271886
rect -7506 264906 -6926 264918
rect 11254 264906 11834 264918
rect 47254 264906 47834 264918
rect 83254 264906 83834 264918
rect 119254 264906 119834 264918
rect 155254 264906 155834 264918
rect 191254 264906 191834 264918
rect 227254 264906 227834 264918
rect 263254 264906 263834 264918
rect 299254 264906 299834 264918
rect 335254 264906 335834 264918
rect 371254 264906 371834 264918
rect 407254 264906 407834 264918
rect 443254 264906 443834 264918
rect 479254 264906 479834 264918
rect 515254 264906 515834 264918
rect 551254 264906 551834 264918
rect 590850 264906 591430 264918
rect -8426 264894 592350 264906
rect -8426 264658 -7334 264894
rect -7098 264658 11426 264894
rect 11662 264658 47426 264894
rect 47662 264658 83426 264894
rect 83662 264658 119426 264894
rect 119662 264658 155426 264894
rect 155662 264658 191426 264894
rect 191662 264658 227426 264894
rect 227662 264658 263426 264894
rect 263662 264658 299426 264894
rect 299662 264658 335426 264894
rect 335662 264658 371426 264894
rect 371662 264658 407426 264894
rect 407662 264658 443426 264894
rect 443662 264658 479426 264894
rect 479662 264658 515426 264894
rect 515662 264658 551426 264894
rect 551662 264658 591022 264894
rect 591258 264658 592350 264894
rect -8426 264574 592350 264658
rect -8426 264338 -7334 264574
rect -7098 264338 11426 264574
rect 11662 264338 47426 264574
rect 47662 264338 83426 264574
rect 83662 264338 119426 264574
rect 119662 264338 155426 264574
rect 155662 264338 191426 264574
rect 191662 264338 227426 264574
rect 227662 264338 263426 264574
rect 263662 264338 299426 264574
rect 299662 264338 335426 264574
rect 335662 264338 371426 264574
rect 371662 264338 407426 264574
rect 407662 264338 443426 264574
rect 443662 264338 479426 264574
rect 479662 264338 515426 264574
rect 515662 264338 551426 264574
rect 551662 264338 591022 264574
rect 591258 264338 592350 264574
rect -8426 264326 592350 264338
rect -7506 264314 -6926 264326
rect 11254 264314 11834 264326
rect 47254 264314 47834 264326
rect 83254 264314 83834 264326
rect 119254 264314 119834 264326
rect 155254 264314 155834 264326
rect 191254 264314 191834 264326
rect 227254 264314 227834 264326
rect 263254 264314 263834 264326
rect 299254 264314 299834 264326
rect 335254 264314 335834 264326
rect 371254 264314 371834 264326
rect 407254 264314 407834 264326
rect 443254 264314 443834 264326
rect 479254 264314 479834 264326
rect 515254 264314 515834 264326
rect 551254 264314 551834 264326
rect 590850 264314 591430 264326
rect -5666 261426 -5086 261438
rect 7774 261426 8354 261438
rect 43774 261426 44354 261438
rect 79774 261426 80354 261438
rect 115774 261426 116354 261438
rect 151774 261426 152354 261438
rect 187774 261426 188354 261438
rect 223774 261426 224354 261438
rect 259774 261426 260354 261438
rect 295774 261426 296354 261438
rect 331774 261426 332354 261438
rect 367774 261426 368354 261438
rect 403774 261426 404354 261438
rect 439774 261426 440354 261438
rect 475774 261426 476354 261438
rect 511774 261426 512354 261438
rect 547774 261426 548354 261438
rect 589010 261426 589590 261438
rect -6586 261414 590510 261426
rect -6586 261178 -5494 261414
rect -5258 261178 7946 261414
rect 8182 261178 43946 261414
rect 44182 261178 79946 261414
rect 80182 261178 115946 261414
rect 116182 261178 151946 261414
rect 152182 261178 187946 261414
rect 188182 261178 223946 261414
rect 224182 261178 259946 261414
rect 260182 261178 295946 261414
rect 296182 261178 331946 261414
rect 332182 261178 367946 261414
rect 368182 261178 403946 261414
rect 404182 261178 439946 261414
rect 440182 261178 475946 261414
rect 476182 261178 511946 261414
rect 512182 261178 547946 261414
rect 548182 261178 589182 261414
rect 589418 261178 590510 261414
rect -6586 261094 590510 261178
rect -6586 260858 -5494 261094
rect -5258 260858 7946 261094
rect 8182 260858 43946 261094
rect 44182 260858 79946 261094
rect 80182 260858 115946 261094
rect 116182 260858 151946 261094
rect 152182 260858 187946 261094
rect 188182 260858 223946 261094
rect 224182 260858 259946 261094
rect 260182 260858 295946 261094
rect 296182 260858 331946 261094
rect 332182 260858 367946 261094
rect 368182 260858 403946 261094
rect 404182 260858 439946 261094
rect 440182 260858 475946 261094
rect 476182 260858 511946 261094
rect 512182 260858 547946 261094
rect 548182 260858 589182 261094
rect 589418 260858 590510 261094
rect -6586 260846 590510 260858
rect -5666 260834 -5086 260846
rect 7774 260834 8354 260846
rect 43774 260834 44354 260846
rect 79774 260834 80354 260846
rect 115774 260834 116354 260846
rect 151774 260834 152354 260846
rect 187774 260834 188354 260846
rect 223774 260834 224354 260846
rect 259774 260834 260354 260846
rect 295774 260834 296354 260846
rect 331774 260834 332354 260846
rect 367774 260834 368354 260846
rect 403774 260834 404354 260846
rect 439774 260834 440354 260846
rect 475774 260834 476354 260846
rect 511774 260834 512354 260846
rect 547774 260834 548354 260846
rect 589010 260834 589590 260846
rect -3826 257946 -3246 257958
rect 4294 257946 4874 257958
rect 40294 257946 40874 257958
rect 76294 257946 76874 257958
rect 112294 257946 112874 257958
rect 148294 257946 148874 257958
rect 184294 257946 184874 257958
rect 220294 257946 220874 257958
rect 256294 257946 256874 257958
rect 292294 257946 292874 257958
rect 328294 257946 328874 257958
rect 364294 257946 364874 257958
rect 400294 257946 400874 257958
rect 436294 257946 436874 257958
rect 472294 257946 472874 257958
rect 508294 257946 508874 257958
rect 544294 257946 544874 257958
rect 580294 257946 580874 257958
rect 587170 257946 587750 257958
rect -4746 257934 588670 257946
rect -4746 257698 -3654 257934
rect -3418 257698 4466 257934
rect 4702 257698 40466 257934
rect 40702 257698 76466 257934
rect 76702 257698 112466 257934
rect 112702 257698 148466 257934
rect 148702 257698 184466 257934
rect 184702 257698 220466 257934
rect 220702 257698 256466 257934
rect 256702 257698 292466 257934
rect 292702 257698 328466 257934
rect 328702 257698 364466 257934
rect 364702 257698 400466 257934
rect 400702 257698 436466 257934
rect 436702 257698 472466 257934
rect 472702 257698 508466 257934
rect 508702 257698 544466 257934
rect 544702 257698 580466 257934
rect 580702 257698 587342 257934
rect 587578 257698 588670 257934
rect -4746 257614 588670 257698
rect -4746 257378 -3654 257614
rect -3418 257378 4466 257614
rect 4702 257378 40466 257614
rect 40702 257378 76466 257614
rect 76702 257378 112466 257614
rect 112702 257378 148466 257614
rect 148702 257378 184466 257614
rect 184702 257378 220466 257614
rect 220702 257378 256466 257614
rect 256702 257378 292466 257614
rect 292702 257378 328466 257614
rect 328702 257378 364466 257614
rect 364702 257378 400466 257614
rect 400702 257378 436466 257614
rect 436702 257378 472466 257614
rect 472702 257378 508466 257614
rect 508702 257378 544466 257614
rect 544702 257378 580466 257614
rect 580702 257378 587342 257614
rect 587578 257378 588670 257614
rect -4746 257366 588670 257378
rect -3826 257354 -3246 257366
rect 4294 257354 4874 257366
rect 40294 257354 40874 257366
rect 76294 257354 76874 257366
rect 112294 257354 112874 257366
rect 148294 257354 148874 257366
rect 184294 257354 184874 257366
rect 220294 257354 220874 257366
rect 256294 257354 256874 257366
rect 292294 257354 292874 257366
rect 328294 257354 328874 257366
rect 364294 257354 364874 257366
rect 400294 257354 400874 257366
rect 436294 257354 436874 257366
rect 472294 257354 472874 257366
rect 508294 257354 508874 257366
rect 544294 257354 544874 257366
rect 580294 257354 580874 257366
rect 587170 257354 587750 257366
rect -1986 254466 -1406 254478
rect 814 254466 1394 254478
rect 36814 254466 37394 254478
rect 72814 254466 73394 254478
rect 108814 254466 109394 254478
rect 144814 254466 145394 254478
rect 180814 254466 181394 254478
rect 216814 254466 217394 254478
rect 252814 254466 253394 254478
rect 288814 254466 289394 254478
rect 324814 254466 325394 254478
rect 360814 254466 361394 254478
rect 396814 254466 397394 254478
rect 432814 254466 433394 254478
rect 468814 254466 469394 254478
rect 504814 254466 505394 254478
rect 540814 254466 541394 254478
rect 576814 254466 577394 254478
rect 585330 254466 585910 254478
rect -2906 254454 586830 254466
rect -2906 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586830 254454
rect -2906 254134 586830 254218
rect -2906 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586830 254134
rect -2906 253886 586830 253898
rect -1986 253874 -1406 253886
rect 814 253874 1394 253886
rect 36814 253874 37394 253886
rect 72814 253874 73394 253886
rect 108814 253874 109394 253886
rect 144814 253874 145394 253886
rect 180814 253874 181394 253886
rect 216814 253874 217394 253886
rect 252814 253874 253394 253886
rect 288814 253874 289394 253886
rect 324814 253874 325394 253886
rect 360814 253874 361394 253886
rect 396814 253874 397394 253886
rect 432814 253874 433394 253886
rect 468814 253874 469394 253886
rect 504814 253874 505394 253886
rect 540814 253874 541394 253886
rect 576814 253874 577394 253886
rect 585330 253874 585910 253886
rect -8426 246906 -7846 246918
rect 29254 246906 29834 246918
rect 65254 246906 65834 246918
rect 101254 246906 101834 246918
rect 137254 246906 137834 246918
rect 173254 246906 173834 246918
rect 209254 246906 209834 246918
rect 245254 246906 245834 246918
rect 281254 246906 281834 246918
rect 317254 246906 317834 246918
rect 353254 246906 353834 246918
rect 389254 246906 389834 246918
rect 425254 246906 425834 246918
rect 461254 246906 461834 246918
rect 497254 246906 497834 246918
rect 533254 246906 533834 246918
rect 569254 246906 569834 246918
rect 591770 246906 592350 246918
rect -8426 246894 592350 246906
rect -8426 246658 -8254 246894
rect -8018 246658 29426 246894
rect 29662 246658 65426 246894
rect 65662 246658 101426 246894
rect 101662 246658 137426 246894
rect 137662 246658 173426 246894
rect 173662 246658 209426 246894
rect 209662 246658 245426 246894
rect 245662 246658 281426 246894
rect 281662 246658 317426 246894
rect 317662 246658 353426 246894
rect 353662 246658 389426 246894
rect 389662 246658 425426 246894
rect 425662 246658 461426 246894
rect 461662 246658 497426 246894
rect 497662 246658 533426 246894
rect 533662 246658 569426 246894
rect 569662 246658 591942 246894
rect 592178 246658 592350 246894
rect -8426 246574 592350 246658
rect -8426 246338 -8254 246574
rect -8018 246338 29426 246574
rect 29662 246338 65426 246574
rect 65662 246338 101426 246574
rect 101662 246338 137426 246574
rect 137662 246338 173426 246574
rect 173662 246338 209426 246574
rect 209662 246338 245426 246574
rect 245662 246338 281426 246574
rect 281662 246338 317426 246574
rect 317662 246338 353426 246574
rect 353662 246338 389426 246574
rect 389662 246338 425426 246574
rect 425662 246338 461426 246574
rect 461662 246338 497426 246574
rect 497662 246338 533426 246574
rect 533662 246338 569426 246574
rect 569662 246338 591942 246574
rect 592178 246338 592350 246574
rect -8426 246326 592350 246338
rect -8426 246314 -7846 246326
rect 29254 246314 29834 246326
rect 65254 246314 65834 246326
rect 101254 246314 101834 246326
rect 137254 246314 137834 246326
rect 173254 246314 173834 246326
rect 209254 246314 209834 246326
rect 245254 246314 245834 246326
rect 281254 246314 281834 246326
rect 317254 246314 317834 246326
rect 353254 246314 353834 246326
rect 389254 246314 389834 246326
rect 425254 246314 425834 246326
rect 461254 246314 461834 246326
rect 497254 246314 497834 246326
rect 533254 246314 533834 246326
rect 569254 246314 569834 246326
rect 591770 246314 592350 246326
rect -6586 243426 -6006 243438
rect 25774 243426 26354 243438
rect 61774 243426 62354 243438
rect 97774 243426 98354 243438
rect 133774 243426 134354 243438
rect 169774 243426 170354 243438
rect 205774 243426 206354 243438
rect 241774 243426 242354 243438
rect 277774 243426 278354 243438
rect 313774 243426 314354 243438
rect 349774 243426 350354 243438
rect 385774 243426 386354 243438
rect 421774 243426 422354 243438
rect 457774 243426 458354 243438
rect 493774 243426 494354 243438
rect 529774 243426 530354 243438
rect 565774 243426 566354 243438
rect 589930 243426 590510 243438
rect -6586 243414 590510 243426
rect -6586 243178 -6414 243414
rect -6178 243178 25946 243414
rect 26182 243178 61946 243414
rect 62182 243178 97946 243414
rect 98182 243178 133946 243414
rect 134182 243178 169946 243414
rect 170182 243178 205946 243414
rect 206182 243178 241946 243414
rect 242182 243178 277946 243414
rect 278182 243178 313946 243414
rect 314182 243178 349946 243414
rect 350182 243178 385946 243414
rect 386182 243178 421946 243414
rect 422182 243178 457946 243414
rect 458182 243178 493946 243414
rect 494182 243178 529946 243414
rect 530182 243178 565946 243414
rect 566182 243178 590102 243414
rect 590338 243178 590510 243414
rect -6586 243094 590510 243178
rect -6586 242858 -6414 243094
rect -6178 242858 25946 243094
rect 26182 242858 61946 243094
rect 62182 242858 97946 243094
rect 98182 242858 133946 243094
rect 134182 242858 169946 243094
rect 170182 242858 205946 243094
rect 206182 242858 241946 243094
rect 242182 242858 277946 243094
rect 278182 242858 313946 243094
rect 314182 242858 349946 243094
rect 350182 242858 385946 243094
rect 386182 242858 421946 243094
rect 422182 242858 457946 243094
rect 458182 242858 493946 243094
rect 494182 242858 529946 243094
rect 530182 242858 565946 243094
rect 566182 242858 590102 243094
rect 590338 242858 590510 243094
rect -6586 242846 590510 242858
rect -6586 242834 -6006 242846
rect 25774 242834 26354 242846
rect 61774 242834 62354 242846
rect 97774 242834 98354 242846
rect 133774 242834 134354 242846
rect 169774 242834 170354 242846
rect 205774 242834 206354 242846
rect 241774 242834 242354 242846
rect 277774 242834 278354 242846
rect 313774 242834 314354 242846
rect 349774 242834 350354 242846
rect 385774 242834 386354 242846
rect 421774 242834 422354 242846
rect 457774 242834 458354 242846
rect 493774 242834 494354 242846
rect 529774 242834 530354 242846
rect 565774 242834 566354 242846
rect 589930 242834 590510 242846
rect -4746 239946 -4166 239958
rect 22294 239946 22874 239958
rect 58294 239946 58874 239958
rect 94294 239946 94874 239958
rect 130294 239946 130874 239958
rect 166294 239946 166874 239958
rect 202294 239946 202874 239958
rect 238294 239946 238874 239958
rect 274294 239946 274874 239958
rect 310294 239946 310874 239958
rect 346294 239946 346874 239958
rect 382294 239946 382874 239958
rect 418294 239946 418874 239958
rect 454294 239946 454874 239958
rect 490294 239946 490874 239958
rect 526294 239946 526874 239958
rect 562294 239946 562874 239958
rect 588090 239946 588670 239958
rect -4746 239934 588670 239946
rect -4746 239698 -4574 239934
rect -4338 239698 22466 239934
rect 22702 239698 58466 239934
rect 58702 239698 94466 239934
rect 94702 239698 130466 239934
rect 130702 239698 166466 239934
rect 166702 239698 202466 239934
rect 202702 239698 238466 239934
rect 238702 239698 274466 239934
rect 274702 239698 310466 239934
rect 310702 239698 346466 239934
rect 346702 239698 382466 239934
rect 382702 239698 418466 239934
rect 418702 239698 454466 239934
rect 454702 239698 490466 239934
rect 490702 239698 526466 239934
rect 526702 239698 562466 239934
rect 562702 239698 588262 239934
rect 588498 239698 588670 239934
rect -4746 239614 588670 239698
rect -4746 239378 -4574 239614
rect -4338 239378 22466 239614
rect 22702 239378 58466 239614
rect 58702 239378 94466 239614
rect 94702 239378 130466 239614
rect 130702 239378 166466 239614
rect 166702 239378 202466 239614
rect 202702 239378 238466 239614
rect 238702 239378 274466 239614
rect 274702 239378 310466 239614
rect 310702 239378 346466 239614
rect 346702 239378 382466 239614
rect 382702 239378 418466 239614
rect 418702 239378 454466 239614
rect 454702 239378 490466 239614
rect 490702 239378 526466 239614
rect 526702 239378 562466 239614
rect 562702 239378 588262 239614
rect 588498 239378 588670 239614
rect -4746 239366 588670 239378
rect -4746 239354 -4166 239366
rect 22294 239354 22874 239366
rect 58294 239354 58874 239366
rect 94294 239354 94874 239366
rect 130294 239354 130874 239366
rect 166294 239354 166874 239366
rect 202294 239354 202874 239366
rect 238294 239354 238874 239366
rect 274294 239354 274874 239366
rect 310294 239354 310874 239366
rect 346294 239354 346874 239366
rect 382294 239354 382874 239366
rect 418294 239354 418874 239366
rect 454294 239354 454874 239366
rect 490294 239354 490874 239366
rect 526294 239354 526874 239366
rect 562294 239354 562874 239366
rect 588090 239354 588670 239366
rect -2906 236466 -2326 236478
rect 18814 236466 19394 236478
rect 54814 236466 55394 236478
rect 90814 236466 91394 236478
rect 126814 236466 127394 236478
rect 162814 236466 163394 236478
rect 198814 236466 199394 236478
rect 234814 236466 235394 236478
rect 270814 236466 271394 236478
rect 306814 236466 307394 236478
rect 342814 236466 343394 236478
rect 378814 236466 379394 236478
rect 414814 236466 415394 236478
rect 450814 236466 451394 236478
rect 486814 236466 487394 236478
rect 522814 236466 523394 236478
rect 558814 236466 559394 236478
rect 586250 236466 586830 236478
rect -2906 236454 586830 236466
rect -2906 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586830 236454
rect -2906 236134 586830 236218
rect -2906 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586830 236134
rect -2906 235886 586830 235898
rect -2906 235874 -2326 235886
rect 18814 235874 19394 235886
rect 54814 235874 55394 235886
rect 90814 235874 91394 235886
rect 126814 235874 127394 235886
rect 162814 235874 163394 235886
rect 198814 235874 199394 235886
rect 234814 235874 235394 235886
rect 270814 235874 271394 235886
rect 306814 235874 307394 235886
rect 342814 235874 343394 235886
rect 378814 235874 379394 235886
rect 414814 235874 415394 235886
rect 450814 235874 451394 235886
rect 486814 235874 487394 235886
rect 522814 235874 523394 235886
rect 558814 235874 559394 235886
rect 586250 235874 586830 235886
rect -7506 228906 -6926 228918
rect 11254 228906 11834 228918
rect 47254 228906 47834 228918
rect 83254 228906 83834 228918
rect 119254 228906 119834 228918
rect 155254 228906 155834 228918
rect 191254 228906 191834 228918
rect 227254 228906 227834 228918
rect 263254 228906 263834 228918
rect 299254 228906 299834 228918
rect 335254 228906 335834 228918
rect 371254 228906 371834 228918
rect 407254 228906 407834 228918
rect 443254 228906 443834 228918
rect 479254 228906 479834 228918
rect 515254 228906 515834 228918
rect 551254 228906 551834 228918
rect 590850 228906 591430 228918
rect -8426 228894 592350 228906
rect -8426 228658 -7334 228894
rect -7098 228658 11426 228894
rect 11662 228658 47426 228894
rect 47662 228658 83426 228894
rect 83662 228658 119426 228894
rect 119662 228658 155426 228894
rect 155662 228658 191426 228894
rect 191662 228658 227426 228894
rect 227662 228658 263426 228894
rect 263662 228658 299426 228894
rect 299662 228658 335426 228894
rect 335662 228658 371426 228894
rect 371662 228658 407426 228894
rect 407662 228658 443426 228894
rect 443662 228658 479426 228894
rect 479662 228658 515426 228894
rect 515662 228658 551426 228894
rect 551662 228658 591022 228894
rect 591258 228658 592350 228894
rect -8426 228574 592350 228658
rect -8426 228338 -7334 228574
rect -7098 228338 11426 228574
rect 11662 228338 47426 228574
rect 47662 228338 83426 228574
rect 83662 228338 119426 228574
rect 119662 228338 155426 228574
rect 155662 228338 191426 228574
rect 191662 228338 227426 228574
rect 227662 228338 263426 228574
rect 263662 228338 299426 228574
rect 299662 228338 335426 228574
rect 335662 228338 371426 228574
rect 371662 228338 407426 228574
rect 407662 228338 443426 228574
rect 443662 228338 479426 228574
rect 479662 228338 515426 228574
rect 515662 228338 551426 228574
rect 551662 228338 591022 228574
rect 591258 228338 592350 228574
rect -8426 228326 592350 228338
rect -7506 228314 -6926 228326
rect 11254 228314 11834 228326
rect 47254 228314 47834 228326
rect 83254 228314 83834 228326
rect 119254 228314 119834 228326
rect 155254 228314 155834 228326
rect 191254 228314 191834 228326
rect 227254 228314 227834 228326
rect 263254 228314 263834 228326
rect 299254 228314 299834 228326
rect 335254 228314 335834 228326
rect 371254 228314 371834 228326
rect 407254 228314 407834 228326
rect 443254 228314 443834 228326
rect 479254 228314 479834 228326
rect 515254 228314 515834 228326
rect 551254 228314 551834 228326
rect 590850 228314 591430 228326
rect -5666 225426 -5086 225438
rect 7774 225426 8354 225438
rect 43774 225426 44354 225438
rect 79774 225426 80354 225438
rect 115774 225426 116354 225438
rect 151774 225426 152354 225438
rect 187774 225426 188354 225438
rect 223774 225426 224354 225438
rect 259774 225426 260354 225438
rect 295774 225426 296354 225438
rect 331774 225426 332354 225438
rect 367774 225426 368354 225438
rect 403774 225426 404354 225438
rect 439774 225426 440354 225438
rect 475774 225426 476354 225438
rect 511774 225426 512354 225438
rect 547774 225426 548354 225438
rect 589010 225426 589590 225438
rect -6586 225414 590510 225426
rect -6586 225178 -5494 225414
rect -5258 225178 7946 225414
rect 8182 225178 43946 225414
rect 44182 225178 79946 225414
rect 80182 225178 115946 225414
rect 116182 225178 151946 225414
rect 152182 225178 187946 225414
rect 188182 225178 223946 225414
rect 224182 225178 259946 225414
rect 260182 225178 295946 225414
rect 296182 225178 331946 225414
rect 332182 225178 367946 225414
rect 368182 225178 403946 225414
rect 404182 225178 439946 225414
rect 440182 225178 475946 225414
rect 476182 225178 511946 225414
rect 512182 225178 547946 225414
rect 548182 225178 589182 225414
rect 589418 225178 590510 225414
rect -6586 225094 590510 225178
rect -6586 224858 -5494 225094
rect -5258 224858 7946 225094
rect 8182 224858 43946 225094
rect 44182 224858 79946 225094
rect 80182 224858 115946 225094
rect 116182 224858 151946 225094
rect 152182 224858 187946 225094
rect 188182 224858 223946 225094
rect 224182 224858 259946 225094
rect 260182 224858 295946 225094
rect 296182 224858 331946 225094
rect 332182 224858 367946 225094
rect 368182 224858 403946 225094
rect 404182 224858 439946 225094
rect 440182 224858 475946 225094
rect 476182 224858 511946 225094
rect 512182 224858 547946 225094
rect 548182 224858 589182 225094
rect 589418 224858 590510 225094
rect -6586 224846 590510 224858
rect -5666 224834 -5086 224846
rect 7774 224834 8354 224846
rect 43774 224834 44354 224846
rect 79774 224834 80354 224846
rect 115774 224834 116354 224846
rect 151774 224834 152354 224846
rect 187774 224834 188354 224846
rect 223774 224834 224354 224846
rect 259774 224834 260354 224846
rect 295774 224834 296354 224846
rect 331774 224834 332354 224846
rect 367774 224834 368354 224846
rect 403774 224834 404354 224846
rect 439774 224834 440354 224846
rect 475774 224834 476354 224846
rect 511774 224834 512354 224846
rect 547774 224834 548354 224846
rect 589010 224834 589590 224846
rect -3826 221946 -3246 221958
rect 4294 221946 4874 221958
rect 40294 221946 40874 221958
rect 76294 221946 76874 221958
rect 112294 221946 112874 221958
rect 148294 221946 148874 221958
rect 184294 221946 184874 221958
rect 220294 221946 220874 221958
rect 256294 221946 256874 221958
rect 292294 221946 292874 221958
rect 328294 221946 328874 221958
rect 364294 221946 364874 221958
rect 400294 221946 400874 221958
rect 436294 221946 436874 221958
rect 472294 221946 472874 221958
rect 508294 221946 508874 221958
rect 544294 221946 544874 221958
rect 580294 221946 580874 221958
rect 587170 221946 587750 221958
rect -4746 221934 588670 221946
rect -4746 221698 -3654 221934
rect -3418 221698 4466 221934
rect 4702 221698 40466 221934
rect 40702 221698 76466 221934
rect 76702 221698 112466 221934
rect 112702 221698 148466 221934
rect 148702 221698 184466 221934
rect 184702 221698 220466 221934
rect 220702 221698 256466 221934
rect 256702 221698 292466 221934
rect 292702 221698 328466 221934
rect 328702 221698 364466 221934
rect 364702 221698 400466 221934
rect 400702 221698 436466 221934
rect 436702 221698 472466 221934
rect 472702 221698 508466 221934
rect 508702 221698 544466 221934
rect 544702 221698 580466 221934
rect 580702 221698 587342 221934
rect 587578 221698 588670 221934
rect -4746 221614 588670 221698
rect -4746 221378 -3654 221614
rect -3418 221378 4466 221614
rect 4702 221378 40466 221614
rect 40702 221378 76466 221614
rect 76702 221378 112466 221614
rect 112702 221378 148466 221614
rect 148702 221378 184466 221614
rect 184702 221378 220466 221614
rect 220702 221378 256466 221614
rect 256702 221378 292466 221614
rect 292702 221378 328466 221614
rect 328702 221378 364466 221614
rect 364702 221378 400466 221614
rect 400702 221378 436466 221614
rect 436702 221378 472466 221614
rect 472702 221378 508466 221614
rect 508702 221378 544466 221614
rect 544702 221378 580466 221614
rect 580702 221378 587342 221614
rect 587578 221378 588670 221614
rect -4746 221366 588670 221378
rect -3826 221354 -3246 221366
rect 4294 221354 4874 221366
rect 40294 221354 40874 221366
rect 76294 221354 76874 221366
rect 112294 221354 112874 221366
rect 148294 221354 148874 221366
rect 184294 221354 184874 221366
rect 220294 221354 220874 221366
rect 256294 221354 256874 221366
rect 292294 221354 292874 221366
rect 328294 221354 328874 221366
rect 364294 221354 364874 221366
rect 400294 221354 400874 221366
rect 436294 221354 436874 221366
rect 472294 221354 472874 221366
rect 508294 221354 508874 221366
rect 544294 221354 544874 221366
rect 580294 221354 580874 221366
rect 587170 221354 587750 221366
rect -1986 218466 -1406 218478
rect 814 218466 1394 218478
rect 36814 218466 37394 218478
rect 72814 218466 73394 218478
rect 108814 218466 109394 218478
rect 144814 218466 145394 218478
rect 180814 218466 181394 218478
rect 216814 218466 217394 218478
rect 252814 218466 253394 218478
rect 288814 218466 289394 218478
rect 324814 218466 325394 218478
rect 360814 218466 361394 218478
rect 396814 218466 397394 218478
rect 432814 218466 433394 218478
rect 468814 218466 469394 218478
rect 504814 218466 505394 218478
rect 540814 218466 541394 218478
rect 576814 218466 577394 218478
rect 585330 218466 585910 218478
rect -2906 218454 586830 218466
rect -2906 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586830 218454
rect -2906 218134 586830 218218
rect -2906 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586830 218134
rect -2906 217886 586830 217898
rect -1986 217874 -1406 217886
rect 814 217874 1394 217886
rect 36814 217874 37394 217886
rect 72814 217874 73394 217886
rect 108814 217874 109394 217886
rect 144814 217874 145394 217886
rect 180814 217874 181394 217886
rect 216814 217874 217394 217886
rect 252814 217874 253394 217886
rect 288814 217874 289394 217886
rect 324814 217874 325394 217886
rect 360814 217874 361394 217886
rect 396814 217874 397394 217886
rect 432814 217874 433394 217886
rect 468814 217874 469394 217886
rect 504814 217874 505394 217886
rect 540814 217874 541394 217886
rect 576814 217874 577394 217886
rect 585330 217874 585910 217886
rect -8426 210906 -7846 210918
rect 29254 210906 29834 210918
rect 65254 210906 65834 210918
rect 101254 210906 101834 210918
rect 137254 210906 137834 210918
rect 173254 210906 173834 210918
rect 209254 210906 209834 210918
rect 245254 210906 245834 210918
rect 281254 210906 281834 210918
rect 317254 210906 317834 210918
rect 353254 210906 353834 210918
rect 389254 210906 389834 210918
rect 425254 210906 425834 210918
rect 461254 210906 461834 210918
rect 497254 210906 497834 210918
rect 533254 210906 533834 210918
rect 569254 210906 569834 210918
rect 591770 210906 592350 210918
rect -8426 210894 592350 210906
rect -8426 210658 -8254 210894
rect -8018 210658 29426 210894
rect 29662 210658 65426 210894
rect 65662 210658 101426 210894
rect 101662 210658 137426 210894
rect 137662 210658 173426 210894
rect 173662 210658 209426 210894
rect 209662 210658 245426 210894
rect 245662 210658 281426 210894
rect 281662 210658 317426 210894
rect 317662 210658 353426 210894
rect 353662 210658 389426 210894
rect 389662 210658 425426 210894
rect 425662 210658 461426 210894
rect 461662 210658 497426 210894
rect 497662 210658 533426 210894
rect 533662 210658 569426 210894
rect 569662 210658 591942 210894
rect 592178 210658 592350 210894
rect -8426 210574 592350 210658
rect -8426 210338 -8254 210574
rect -8018 210338 29426 210574
rect 29662 210338 65426 210574
rect 65662 210338 101426 210574
rect 101662 210338 137426 210574
rect 137662 210338 173426 210574
rect 173662 210338 209426 210574
rect 209662 210338 245426 210574
rect 245662 210338 281426 210574
rect 281662 210338 317426 210574
rect 317662 210338 353426 210574
rect 353662 210338 389426 210574
rect 389662 210338 425426 210574
rect 425662 210338 461426 210574
rect 461662 210338 497426 210574
rect 497662 210338 533426 210574
rect 533662 210338 569426 210574
rect 569662 210338 591942 210574
rect 592178 210338 592350 210574
rect -8426 210326 592350 210338
rect -8426 210314 -7846 210326
rect 29254 210314 29834 210326
rect 65254 210314 65834 210326
rect 101254 210314 101834 210326
rect 137254 210314 137834 210326
rect 173254 210314 173834 210326
rect 209254 210314 209834 210326
rect 245254 210314 245834 210326
rect 281254 210314 281834 210326
rect 317254 210314 317834 210326
rect 353254 210314 353834 210326
rect 389254 210314 389834 210326
rect 425254 210314 425834 210326
rect 461254 210314 461834 210326
rect 497254 210314 497834 210326
rect 533254 210314 533834 210326
rect 569254 210314 569834 210326
rect 591770 210314 592350 210326
rect -6586 207426 -6006 207438
rect 25774 207426 26354 207438
rect 61774 207426 62354 207438
rect 97774 207426 98354 207438
rect 133774 207426 134354 207438
rect 169774 207426 170354 207438
rect 205774 207426 206354 207438
rect 241774 207426 242354 207438
rect 277774 207426 278354 207438
rect 313774 207426 314354 207438
rect 349774 207426 350354 207438
rect 385774 207426 386354 207438
rect 421774 207426 422354 207438
rect 457774 207426 458354 207438
rect 493774 207426 494354 207438
rect 529774 207426 530354 207438
rect 565774 207426 566354 207438
rect 589930 207426 590510 207438
rect -6586 207414 590510 207426
rect -6586 207178 -6414 207414
rect -6178 207178 25946 207414
rect 26182 207178 61946 207414
rect 62182 207178 97946 207414
rect 98182 207178 133946 207414
rect 134182 207178 169946 207414
rect 170182 207178 205946 207414
rect 206182 207178 241946 207414
rect 242182 207178 277946 207414
rect 278182 207178 313946 207414
rect 314182 207178 349946 207414
rect 350182 207178 385946 207414
rect 386182 207178 421946 207414
rect 422182 207178 457946 207414
rect 458182 207178 493946 207414
rect 494182 207178 529946 207414
rect 530182 207178 565946 207414
rect 566182 207178 590102 207414
rect 590338 207178 590510 207414
rect -6586 207094 590510 207178
rect -6586 206858 -6414 207094
rect -6178 206858 25946 207094
rect 26182 206858 61946 207094
rect 62182 206858 97946 207094
rect 98182 206858 133946 207094
rect 134182 206858 169946 207094
rect 170182 206858 205946 207094
rect 206182 206858 241946 207094
rect 242182 206858 277946 207094
rect 278182 206858 313946 207094
rect 314182 206858 349946 207094
rect 350182 206858 385946 207094
rect 386182 206858 421946 207094
rect 422182 206858 457946 207094
rect 458182 206858 493946 207094
rect 494182 206858 529946 207094
rect 530182 206858 565946 207094
rect 566182 206858 590102 207094
rect 590338 206858 590510 207094
rect -6586 206846 590510 206858
rect -6586 206834 -6006 206846
rect 25774 206834 26354 206846
rect 61774 206834 62354 206846
rect 97774 206834 98354 206846
rect 133774 206834 134354 206846
rect 169774 206834 170354 206846
rect 205774 206834 206354 206846
rect 241774 206834 242354 206846
rect 277774 206834 278354 206846
rect 313774 206834 314354 206846
rect 349774 206834 350354 206846
rect 385774 206834 386354 206846
rect 421774 206834 422354 206846
rect 457774 206834 458354 206846
rect 493774 206834 494354 206846
rect 529774 206834 530354 206846
rect 565774 206834 566354 206846
rect 589930 206834 590510 206846
rect -4746 203946 -4166 203958
rect 22294 203946 22874 203958
rect 58294 203946 58874 203958
rect 94294 203946 94874 203958
rect 130294 203946 130874 203958
rect 166294 203946 166874 203958
rect 202294 203946 202874 203958
rect 238294 203946 238874 203958
rect 274294 203946 274874 203958
rect 310294 203946 310874 203958
rect 346294 203946 346874 203958
rect 382294 203946 382874 203958
rect 418294 203946 418874 203958
rect 454294 203946 454874 203958
rect 490294 203946 490874 203958
rect 526294 203946 526874 203958
rect 562294 203946 562874 203958
rect 588090 203946 588670 203958
rect -4746 203934 588670 203946
rect -4746 203698 -4574 203934
rect -4338 203698 22466 203934
rect 22702 203698 58466 203934
rect 58702 203698 94466 203934
rect 94702 203698 130466 203934
rect 130702 203698 166466 203934
rect 166702 203698 202466 203934
rect 202702 203698 238466 203934
rect 238702 203698 274466 203934
rect 274702 203698 310466 203934
rect 310702 203698 346466 203934
rect 346702 203698 382466 203934
rect 382702 203698 418466 203934
rect 418702 203698 454466 203934
rect 454702 203698 490466 203934
rect 490702 203698 526466 203934
rect 526702 203698 562466 203934
rect 562702 203698 588262 203934
rect 588498 203698 588670 203934
rect -4746 203614 588670 203698
rect -4746 203378 -4574 203614
rect -4338 203378 22466 203614
rect 22702 203378 58466 203614
rect 58702 203378 94466 203614
rect 94702 203378 130466 203614
rect 130702 203378 166466 203614
rect 166702 203378 202466 203614
rect 202702 203378 238466 203614
rect 238702 203378 274466 203614
rect 274702 203378 310466 203614
rect 310702 203378 346466 203614
rect 346702 203378 382466 203614
rect 382702 203378 418466 203614
rect 418702 203378 454466 203614
rect 454702 203378 490466 203614
rect 490702 203378 526466 203614
rect 526702 203378 562466 203614
rect 562702 203378 588262 203614
rect 588498 203378 588670 203614
rect -4746 203366 588670 203378
rect -4746 203354 -4166 203366
rect 22294 203354 22874 203366
rect 58294 203354 58874 203366
rect 94294 203354 94874 203366
rect 130294 203354 130874 203366
rect 166294 203354 166874 203366
rect 202294 203354 202874 203366
rect 238294 203354 238874 203366
rect 274294 203354 274874 203366
rect 310294 203354 310874 203366
rect 346294 203354 346874 203366
rect 382294 203354 382874 203366
rect 418294 203354 418874 203366
rect 454294 203354 454874 203366
rect 490294 203354 490874 203366
rect 526294 203354 526874 203366
rect 562294 203354 562874 203366
rect 588090 203354 588670 203366
rect -2906 200466 -2326 200478
rect 18814 200466 19394 200478
rect 54814 200466 55394 200478
rect 90814 200466 91394 200478
rect 126814 200466 127394 200478
rect 162814 200466 163394 200478
rect 198814 200466 199394 200478
rect 234814 200466 235394 200478
rect 270814 200466 271394 200478
rect 306814 200466 307394 200478
rect 342814 200466 343394 200478
rect 378814 200466 379394 200478
rect 414814 200466 415394 200478
rect 450814 200466 451394 200478
rect 486814 200466 487394 200478
rect 522814 200466 523394 200478
rect 558814 200466 559394 200478
rect 586250 200466 586830 200478
rect -2906 200454 586830 200466
rect -2906 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586830 200454
rect -2906 200134 586830 200218
rect -2906 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586830 200134
rect -2906 199886 586830 199898
rect -2906 199874 -2326 199886
rect 18814 199874 19394 199886
rect 54814 199874 55394 199886
rect 90814 199874 91394 199886
rect 126814 199874 127394 199886
rect 162814 199874 163394 199886
rect 198814 199874 199394 199886
rect 234814 199874 235394 199886
rect 270814 199874 271394 199886
rect 306814 199874 307394 199886
rect 342814 199874 343394 199886
rect 378814 199874 379394 199886
rect 414814 199874 415394 199886
rect 450814 199874 451394 199886
rect 486814 199874 487394 199886
rect 522814 199874 523394 199886
rect 558814 199874 559394 199886
rect 586250 199874 586830 199886
rect -7506 192906 -6926 192918
rect 11254 192906 11834 192918
rect 47254 192906 47834 192918
rect 83254 192906 83834 192918
rect 119254 192906 119834 192918
rect 155254 192906 155834 192918
rect 191254 192906 191834 192918
rect 227254 192906 227834 192918
rect 263254 192906 263834 192918
rect 299254 192906 299834 192918
rect 335254 192906 335834 192918
rect 371254 192906 371834 192918
rect 407254 192906 407834 192918
rect 443254 192906 443834 192918
rect 479254 192906 479834 192918
rect 515254 192906 515834 192918
rect 551254 192906 551834 192918
rect 590850 192906 591430 192918
rect -8426 192894 592350 192906
rect -8426 192658 -7334 192894
rect -7098 192658 11426 192894
rect 11662 192658 47426 192894
rect 47662 192658 83426 192894
rect 83662 192658 119426 192894
rect 119662 192658 155426 192894
rect 155662 192658 191426 192894
rect 191662 192658 227426 192894
rect 227662 192658 263426 192894
rect 263662 192658 299426 192894
rect 299662 192658 335426 192894
rect 335662 192658 371426 192894
rect 371662 192658 407426 192894
rect 407662 192658 443426 192894
rect 443662 192658 479426 192894
rect 479662 192658 515426 192894
rect 515662 192658 551426 192894
rect 551662 192658 591022 192894
rect 591258 192658 592350 192894
rect -8426 192574 592350 192658
rect -8426 192338 -7334 192574
rect -7098 192338 11426 192574
rect 11662 192338 47426 192574
rect 47662 192338 83426 192574
rect 83662 192338 119426 192574
rect 119662 192338 155426 192574
rect 155662 192338 191426 192574
rect 191662 192338 227426 192574
rect 227662 192338 263426 192574
rect 263662 192338 299426 192574
rect 299662 192338 335426 192574
rect 335662 192338 371426 192574
rect 371662 192338 407426 192574
rect 407662 192338 443426 192574
rect 443662 192338 479426 192574
rect 479662 192338 515426 192574
rect 515662 192338 551426 192574
rect 551662 192338 591022 192574
rect 591258 192338 592350 192574
rect -8426 192326 592350 192338
rect -7506 192314 -6926 192326
rect 11254 192314 11834 192326
rect 47254 192314 47834 192326
rect 83254 192314 83834 192326
rect 119254 192314 119834 192326
rect 155254 192314 155834 192326
rect 191254 192314 191834 192326
rect 227254 192314 227834 192326
rect 263254 192314 263834 192326
rect 299254 192314 299834 192326
rect 335254 192314 335834 192326
rect 371254 192314 371834 192326
rect 407254 192314 407834 192326
rect 443254 192314 443834 192326
rect 479254 192314 479834 192326
rect 515254 192314 515834 192326
rect 551254 192314 551834 192326
rect 590850 192314 591430 192326
rect -5666 189426 -5086 189438
rect 7774 189426 8354 189438
rect 43774 189426 44354 189438
rect 79774 189426 80354 189438
rect 115774 189426 116354 189438
rect 151774 189426 152354 189438
rect 187774 189426 188354 189438
rect 223774 189426 224354 189438
rect 259774 189426 260354 189438
rect 295774 189426 296354 189438
rect 331774 189426 332354 189438
rect 367774 189426 368354 189438
rect 403774 189426 404354 189438
rect 439774 189426 440354 189438
rect 475774 189426 476354 189438
rect 511774 189426 512354 189438
rect 547774 189426 548354 189438
rect 589010 189426 589590 189438
rect -6586 189414 590510 189426
rect -6586 189178 -5494 189414
rect -5258 189178 7946 189414
rect 8182 189178 43946 189414
rect 44182 189178 79946 189414
rect 80182 189178 115946 189414
rect 116182 189178 151946 189414
rect 152182 189178 187946 189414
rect 188182 189178 223946 189414
rect 224182 189178 259946 189414
rect 260182 189178 295946 189414
rect 296182 189178 331946 189414
rect 332182 189178 367946 189414
rect 368182 189178 403946 189414
rect 404182 189178 439946 189414
rect 440182 189178 475946 189414
rect 476182 189178 511946 189414
rect 512182 189178 547946 189414
rect 548182 189178 589182 189414
rect 589418 189178 590510 189414
rect -6586 189094 590510 189178
rect -6586 188858 -5494 189094
rect -5258 188858 7946 189094
rect 8182 188858 43946 189094
rect 44182 188858 79946 189094
rect 80182 188858 115946 189094
rect 116182 188858 151946 189094
rect 152182 188858 187946 189094
rect 188182 188858 223946 189094
rect 224182 188858 259946 189094
rect 260182 188858 295946 189094
rect 296182 188858 331946 189094
rect 332182 188858 367946 189094
rect 368182 188858 403946 189094
rect 404182 188858 439946 189094
rect 440182 188858 475946 189094
rect 476182 188858 511946 189094
rect 512182 188858 547946 189094
rect 548182 188858 589182 189094
rect 589418 188858 590510 189094
rect -6586 188846 590510 188858
rect -5666 188834 -5086 188846
rect 7774 188834 8354 188846
rect 43774 188834 44354 188846
rect 79774 188834 80354 188846
rect 115774 188834 116354 188846
rect 151774 188834 152354 188846
rect 187774 188834 188354 188846
rect 223774 188834 224354 188846
rect 259774 188834 260354 188846
rect 295774 188834 296354 188846
rect 331774 188834 332354 188846
rect 367774 188834 368354 188846
rect 403774 188834 404354 188846
rect 439774 188834 440354 188846
rect 475774 188834 476354 188846
rect 511774 188834 512354 188846
rect 547774 188834 548354 188846
rect 589010 188834 589590 188846
rect -3826 185946 -3246 185958
rect 4294 185946 4874 185958
rect 40294 185946 40874 185958
rect 76294 185946 76874 185958
rect 112294 185946 112874 185958
rect 148294 185946 148874 185958
rect 184294 185946 184874 185958
rect 220294 185946 220874 185958
rect 256294 185946 256874 185958
rect 292294 185946 292874 185958
rect 328294 185946 328874 185958
rect 364294 185946 364874 185958
rect 400294 185946 400874 185958
rect 436294 185946 436874 185958
rect 472294 185946 472874 185958
rect 508294 185946 508874 185958
rect 544294 185946 544874 185958
rect 580294 185946 580874 185958
rect 587170 185946 587750 185958
rect -4746 185934 588670 185946
rect -4746 185698 -3654 185934
rect -3418 185698 4466 185934
rect 4702 185698 40466 185934
rect 40702 185698 76466 185934
rect 76702 185698 112466 185934
rect 112702 185698 148466 185934
rect 148702 185698 184466 185934
rect 184702 185698 220466 185934
rect 220702 185698 256466 185934
rect 256702 185698 292466 185934
rect 292702 185698 328466 185934
rect 328702 185698 364466 185934
rect 364702 185698 400466 185934
rect 400702 185698 436466 185934
rect 436702 185698 472466 185934
rect 472702 185698 508466 185934
rect 508702 185698 544466 185934
rect 544702 185698 580466 185934
rect 580702 185698 587342 185934
rect 587578 185698 588670 185934
rect -4746 185614 588670 185698
rect -4746 185378 -3654 185614
rect -3418 185378 4466 185614
rect 4702 185378 40466 185614
rect 40702 185378 76466 185614
rect 76702 185378 112466 185614
rect 112702 185378 148466 185614
rect 148702 185378 184466 185614
rect 184702 185378 220466 185614
rect 220702 185378 256466 185614
rect 256702 185378 292466 185614
rect 292702 185378 328466 185614
rect 328702 185378 364466 185614
rect 364702 185378 400466 185614
rect 400702 185378 436466 185614
rect 436702 185378 472466 185614
rect 472702 185378 508466 185614
rect 508702 185378 544466 185614
rect 544702 185378 580466 185614
rect 580702 185378 587342 185614
rect 587578 185378 588670 185614
rect -4746 185366 588670 185378
rect -3826 185354 -3246 185366
rect 4294 185354 4874 185366
rect 40294 185354 40874 185366
rect 76294 185354 76874 185366
rect 112294 185354 112874 185366
rect 148294 185354 148874 185366
rect 184294 185354 184874 185366
rect 220294 185354 220874 185366
rect 256294 185354 256874 185366
rect 292294 185354 292874 185366
rect 328294 185354 328874 185366
rect 364294 185354 364874 185366
rect 400294 185354 400874 185366
rect 436294 185354 436874 185366
rect 472294 185354 472874 185366
rect 508294 185354 508874 185366
rect 544294 185354 544874 185366
rect 580294 185354 580874 185366
rect 587170 185354 587750 185366
rect -1986 182466 -1406 182478
rect 814 182466 1394 182478
rect 36814 182466 37394 182478
rect 72814 182466 73394 182478
rect 108814 182466 109394 182478
rect 144814 182466 145394 182478
rect 180814 182466 181394 182478
rect 216814 182466 217394 182478
rect 252814 182466 253394 182478
rect 288814 182466 289394 182478
rect 324814 182466 325394 182478
rect 360814 182466 361394 182478
rect 396814 182466 397394 182478
rect 432814 182466 433394 182478
rect 468814 182466 469394 182478
rect 504814 182466 505394 182478
rect 540814 182466 541394 182478
rect 576814 182466 577394 182478
rect 585330 182466 585910 182478
rect -2906 182454 586830 182466
rect -2906 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586830 182454
rect -2906 182134 586830 182218
rect -2906 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586830 182134
rect -2906 181886 586830 181898
rect -1986 181874 -1406 181886
rect 814 181874 1394 181886
rect 36814 181874 37394 181886
rect 72814 181874 73394 181886
rect 108814 181874 109394 181886
rect 144814 181874 145394 181886
rect 180814 181874 181394 181886
rect 216814 181874 217394 181886
rect 252814 181874 253394 181886
rect 288814 181874 289394 181886
rect 324814 181874 325394 181886
rect 360814 181874 361394 181886
rect 396814 181874 397394 181886
rect 432814 181874 433394 181886
rect 468814 181874 469394 181886
rect 504814 181874 505394 181886
rect 540814 181874 541394 181886
rect 576814 181874 577394 181886
rect 585330 181874 585910 181886
rect -8426 174906 -7846 174918
rect 29254 174906 29834 174918
rect 65254 174906 65834 174918
rect 101254 174906 101834 174918
rect 137254 174906 137834 174918
rect 173254 174906 173834 174918
rect 209254 174906 209834 174918
rect 245254 174906 245834 174918
rect 281254 174906 281834 174918
rect 317254 174906 317834 174918
rect 353254 174906 353834 174918
rect 389254 174906 389834 174918
rect 425254 174906 425834 174918
rect 461254 174906 461834 174918
rect 497254 174906 497834 174918
rect 533254 174906 533834 174918
rect 569254 174906 569834 174918
rect 591770 174906 592350 174918
rect -8426 174894 592350 174906
rect -8426 174658 -8254 174894
rect -8018 174658 29426 174894
rect 29662 174658 65426 174894
rect 65662 174658 101426 174894
rect 101662 174658 137426 174894
rect 137662 174658 173426 174894
rect 173662 174658 209426 174894
rect 209662 174658 245426 174894
rect 245662 174658 281426 174894
rect 281662 174658 317426 174894
rect 317662 174658 353426 174894
rect 353662 174658 389426 174894
rect 389662 174658 425426 174894
rect 425662 174658 461426 174894
rect 461662 174658 497426 174894
rect 497662 174658 533426 174894
rect 533662 174658 569426 174894
rect 569662 174658 591942 174894
rect 592178 174658 592350 174894
rect -8426 174574 592350 174658
rect -8426 174338 -8254 174574
rect -8018 174338 29426 174574
rect 29662 174338 65426 174574
rect 65662 174338 101426 174574
rect 101662 174338 137426 174574
rect 137662 174338 173426 174574
rect 173662 174338 209426 174574
rect 209662 174338 245426 174574
rect 245662 174338 281426 174574
rect 281662 174338 317426 174574
rect 317662 174338 353426 174574
rect 353662 174338 389426 174574
rect 389662 174338 425426 174574
rect 425662 174338 461426 174574
rect 461662 174338 497426 174574
rect 497662 174338 533426 174574
rect 533662 174338 569426 174574
rect 569662 174338 591942 174574
rect 592178 174338 592350 174574
rect -8426 174326 592350 174338
rect -8426 174314 -7846 174326
rect 29254 174314 29834 174326
rect 65254 174314 65834 174326
rect 101254 174314 101834 174326
rect 137254 174314 137834 174326
rect 173254 174314 173834 174326
rect 209254 174314 209834 174326
rect 245254 174314 245834 174326
rect 281254 174314 281834 174326
rect 317254 174314 317834 174326
rect 353254 174314 353834 174326
rect 389254 174314 389834 174326
rect 425254 174314 425834 174326
rect 461254 174314 461834 174326
rect 497254 174314 497834 174326
rect 533254 174314 533834 174326
rect 569254 174314 569834 174326
rect 591770 174314 592350 174326
rect -6586 171426 -6006 171438
rect 25774 171426 26354 171438
rect 61774 171426 62354 171438
rect 97774 171426 98354 171438
rect 133774 171426 134354 171438
rect 169774 171426 170354 171438
rect 205774 171426 206354 171438
rect 241774 171426 242354 171438
rect 277774 171426 278354 171438
rect 313774 171426 314354 171438
rect 349774 171426 350354 171438
rect 385774 171426 386354 171438
rect 421774 171426 422354 171438
rect 457774 171426 458354 171438
rect 493774 171426 494354 171438
rect 529774 171426 530354 171438
rect 565774 171426 566354 171438
rect 589930 171426 590510 171438
rect -6586 171414 590510 171426
rect -6586 171178 -6414 171414
rect -6178 171178 25946 171414
rect 26182 171178 61946 171414
rect 62182 171178 97946 171414
rect 98182 171178 133946 171414
rect 134182 171178 169946 171414
rect 170182 171178 205946 171414
rect 206182 171178 241946 171414
rect 242182 171178 277946 171414
rect 278182 171178 313946 171414
rect 314182 171178 349946 171414
rect 350182 171178 385946 171414
rect 386182 171178 421946 171414
rect 422182 171178 457946 171414
rect 458182 171178 493946 171414
rect 494182 171178 529946 171414
rect 530182 171178 565946 171414
rect 566182 171178 590102 171414
rect 590338 171178 590510 171414
rect -6586 171094 590510 171178
rect -6586 170858 -6414 171094
rect -6178 170858 25946 171094
rect 26182 170858 61946 171094
rect 62182 170858 97946 171094
rect 98182 170858 133946 171094
rect 134182 170858 169946 171094
rect 170182 170858 205946 171094
rect 206182 170858 241946 171094
rect 242182 170858 277946 171094
rect 278182 170858 313946 171094
rect 314182 170858 349946 171094
rect 350182 170858 385946 171094
rect 386182 170858 421946 171094
rect 422182 170858 457946 171094
rect 458182 170858 493946 171094
rect 494182 170858 529946 171094
rect 530182 170858 565946 171094
rect 566182 170858 590102 171094
rect 590338 170858 590510 171094
rect -6586 170846 590510 170858
rect -6586 170834 -6006 170846
rect 25774 170834 26354 170846
rect 61774 170834 62354 170846
rect 97774 170834 98354 170846
rect 133774 170834 134354 170846
rect 169774 170834 170354 170846
rect 205774 170834 206354 170846
rect 241774 170834 242354 170846
rect 277774 170834 278354 170846
rect 313774 170834 314354 170846
rect 349774 170834 350354 170846
rect 385774 170834 386354 170846
rect 421774 170834 422354 170846
rect 457774 170834 458354 170846
rect 493774 170834 494354 170846
rect 529774 170834 530354 170846
rect 565774 170834 566354 170846
rect 589930 170834 590510 170846
rect -4746 167946 -4166 167958
rect 22294 167946 22874 167958
rect 58294 167946 58874 167958
rect 94294 167946 94874 167958
rect 130294 167946 130874 167958
rect 166294 167946 166874 167958
rect 202294 167946 202874 167958
rect 238294 167946 238874 167958
rect 274294 167946 274874 167958
rect 310294 167946 310874 167958
rect 346294 167946 346874 167958
rect 382294 167946 382874 167958
rect 418294 167946 418874 167958
rect 454294 167946 454874 167958
rect 490294 167946 490874 167958
rect 526294 167946 526874 167958
rect 562294 167946 562874 167958
rect 588090 167946 588670 167958
rect -4746 167934 588670 167946
rect -4746 167698 -4574 167934
rect -4338 167698 22466 167934
rect 22702 167698 58466 167934
rect 58702 167698 94466 167934
rect 94702 167698 130466 167934
rect 130702 167698 166466 167934
rect 166702 167698 202466 167934
rect 202702 167698 238466 167934
rect 238702 167698 274466 167934
rect 274702 167698 310466 167934
rect 310702 167698 346466 167934
rect 346702 167698 382466 167934
rect 382702 167698 418466 167934
rect 418702 167698 454466 167934
rect 454702 167698 490466 167934
rect 490702 167698 526466 167934
rect 526702 167698 562466 167934
rect 562702 167698 588262 167934
rect 588498 167698 588670 167934
rect -4746 167614 588670 167698
rect -4746 167378 -4574 167614
rect -4338 167378 22466 167614
rect 22702 167378 58466 167614
rect 58702 167378 94466 167614
rect 94702 167378 130466 167614
rect 130702 167378 166466 167614
rect 166702 167378 202466 167614
rect 202702 167378 238466 167614
rect 238702 167378 274466 167614
rect 274702 167378 310466 167614
rect 310702 167378 346466 167614
rect 346702 167378 382466 167614
rect 382702 167378 418466 167614
rect 418702 167378 454466 167614
rect 454702 167378 490466 167614
rect 490702 167378 526466 167614
rect 526702 167378 562466 167614
rect 562702 167378 588262 167614
rect 588498 167378 588670 167614
rect -4746 167366 588670 167378
rect -4746 167354 -4166 167366
rect 22294 167354 22874 167366
rect 58294 167354 58874 167366
rect 94294 167354 94874 167366
rect 130294 167354 130874 167366
rect 166294 167354 166874 167366
rect 202294 167354 202874 167366
rect 238294 167354 238874 167366
rect 274294 167354 274874 167366
rect 310294 167354 310874 167366
rect 346294 167354 346874 167366
rect 382294 167354 382874 167366
rect 418294 167354 418874 167366
rect 454294 167354 454874 167366
rect 490294 167354 490874 167366
rect 526294 167354 526874 167366
rect 562294 167354 562874 167366
rect 588090 167354 588670 167366
rect -2906 164466 -2326 164478
rect 18814 164466 19394 164478
rect 54814 164466 55394 164478
rect 90814 164466 91394 164478
rect 126814 164466 127394 164478
rect 162814 164466 163394 164478
rect 198814 164466 199394 164478
rect 234814 164466 235394 164478
rect 270814 164466 271394 164478
rect 306814 164466 307394 164478
rect 342814 164466 343394 164478
rect 378814 164466 379394 164478
rect 414814 164466 415394 164478
rect 450814 164466 451394 164478
rect 486814 164466 487394 164478
rect 522814 164466 523394 164478
rect 558814 164466 559394 164478
rect 586250 164466 586830 164478
rect -2906 164454 586830 164466
rect -2906 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586830 164454
rect -2906 164134 586830 164218
rect -2906 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586830 164134
rect -2906 163886 586830 163898
rect -2906 163874 -2326 163886
rect 18814 163874 19394 163886
rect 54814 163874 55394 163886
rect 90814 163874 91394 163886
rect 126814 163874 127394 163886
rect 162814 163874 163394 163886
rect 198814 163874 199394 163886
rect 234814 163874 235394 163886
rect 270814 163874 271394 163886
rect 306814 163874 307394 163886
rect 342814 163874 343394 163886
rect 378814 163874 379394 163886
rect 414814 163874 415394 163886
rect 450814 163874 451394 163886
rect 486814 163874 487394 163886
rect 522814 163874 523394 163886
rect 558814 163874 559394 163886
rect 586250 163874 586830 163886
rect -7506 156906 -6926 156918
rect 11254 156906 11834 156918
rect 47254 156906 47834 156918
rect 83254 156906 83834 156918
rect 119254 156906 119834 156918
rect 155254 156906 155834 156918
rect 191254 156906 191834 156918
rect 227254 156906 227834 156918
rect 263254 156906 263834 156918
rect 299254 156906 299834 156918
rect 335254 156906 335834 156918
rect 371254 156906 371834 156918
rect 407254 156906 407834 156918
rect 443254 156906 443834 156918
rect 479254 156906 479834 156918
rect 515254 156906 515834 156918
rect 551254 156906 551834 156918
rect 590850 156906 591430 156918
rect -8426 156894 592350 156906
rect -8426 156658 -7334 156894
rect -7098 156658 11426 156894
rect 11662 156658 47426 156894
rect 47662 156658 83426 156894
rect 83662 156658 119426 156894
rect 119662 156658 155426 156894
rect 155662 156658 191426 156894
rect 191662 156658 227426 156894
rect 227662 156658 263426 156894
rect 263662 156658 299426 156894
rect 299662 156658 335426 156894
rect 335662 156658 371426 156894
rect 371662 156658 407426 156894
rect 407662 156658 443426 156894
rect 443662 156658 479426 156894
rect 479662 156658 515426 156894
rect 515662 156658 551426 156894
rect 551662 156658 591022 156894
rect 591258 156658 592350 156894
rect -8426 156574 592350 156658
rect -8426 156338 -7334 156574
rect -7098 156338 11426 156574
rect 11662 156338 47426 156574
rect 47662 156338 83426 156574
rect 83662 156338 119426 156574
rect 119662 156338 155426 156574
rect 155662 156338 191426 156574
rect 191662 156338 227426 156574
rect 227662 156338 263426 156574
rect 263662 156338 299426 156574
rect 299662 156338 335426 156574
rect 335662 156338 371426 156574
rect 371662 156338 407426 156574
rect 407662 156338 443426 156574
rect 443662 156338 479426 156574
rect 479662 156338 515426 156574
rect 515662 156338 551426 156574
rect 551662 156338 591022 156574
rect 591258 156338 592350 156574
rect -8426 156326 592350 156338
rect -7506 156314 -6926 156326
rect 11254 156314 11834 156326
rect 47254 156314 47834 156326
rect 83254 156314 83834 156326
rect 119254 156314 119834 156326
rect 155254 156314 155834 156326
rect 191254 156314 191834 156326
rect 227254 156314 227834 156326
rect 263254 156314 263834 156326
rect 299254 156314 299834 156326
rect 335254 156314 335834 156326
rect 371254 156314 371834 156326
rect 407254 156314 407834 156326
rect 443254 156314 443834 156326
rect 479254 156314 479834 156326
rect 515254 156314 515834 156326
rect 551254 156314 551834 156326
rect 590850 156314 591430 156326
rect -5666 153426 -5086 153438
rect 7774 153426 8354 153438
rect 43774 153426 44354 153438
rect 79774 153426 80354 153438
rect 115774 153426 116354 153438
rect 151774 153426 152354 153438
rect 187774 153426 188354 153438
rect 223774 153426 224354 153438
rect 259774 153426 260354 153438
rect 295774 153426 296354 153438
rect 331774 153426 332354 153438
rect 367774 153426 368354 153438
rect 403774 153426 404354 153438
rect 439774 153426 440354 153438
rect 475774 153426 476354 153438
rect 511774 153426 512354 153438
rect 547774 153426 548354 153438
rect 589010 153426 589590 153438
rect -6586 153414 590510 153426
rect -6586 153178 -5494 153414
rect -5258 153178 7946 153414
rect 8182 153178 43946 153414
rect 44182 153178 79946 153414
rect 80182 153178 115946 153414
rect 116182 153178 151946 153414
rect 152182 153178 187946 153414
rect 188182 153178 223946 153414
rect 224182 153178 259946 153414
rect 260182 153178 295946 153414
rect 296182 153178 331946 153414
rect 332182 153178 367946 153414
rect 368182 153178 403946 153414
rect 404182 153178 439946 153414
rect 440182 153178 475946 153414
rect 476182 153178 511946 153414
rect 512182 153178 547946 153414
rect 548182 153178 589182 153414
rect 589418 153178 590510 153414
rect -6586 153094 590510 153178
rect -6586 152858 -5494 153094
rect -5258 152858 7946 153094
rect 8182 152858 43946 153094
rect 44182 152858 79946 153094
rect 80182 152858 115946 153094
rect 116182 152858 151946 153094
rect 152182 152858 187946 153094
rect 188182 152858 223946 153094
rect 224182 152858 259946 153094
rect 260182 152858 295946 153094
rect 296182 152858 331946 153094
rect 332182 152858 367946 153094
rect 368182 152858 403946 153094
rect 404182 152858 439946 153094
rect 440182 152858 475946 153094
rect 476182 152858 511946 153094
rect 512182 152858 547946 153094
rect 548182 152858 589182 153094
rect 589418 152858 590510 153094
rect -6586 152846 590510 152858
rect -5666 152834 -5086 152846
rect 7774 152834 8354 152846
rect 43774 152834 44354 152846
rect 79774 152834 80354 152846
rect 115774 152834 116354 152846
rect 151774 152834 152354 152846
rect 187774 152834 188354 152846
rect 223774 152834 224354 152846
rect 259774 152834 260354 152846
rect 295774 152834 296354 152846
rect 331774 152834 332354 152846
rect 367774 152834 368354 152846
rect 403774 152834 404354 152846
rect 439774 152834 440354 152846
rect 475774 152834 476354 152846
rect 511774 152834 512354 152846
rect 547774 152834 548354 152846
rect 589010 152834 589590 152846
rect -3826 149946 -3246 149958
rect 4294 149946 4874 149958
rect 40294 149946 40874 149958
rect 76294 149946 76874 149958
rect 112294 149946 112874 149958
rect 148294 149946 148874 149958
rect 184294 149946 184874 149958
rect 220294 149946 220874 149958
rect 256294 149946 256874 149958
rect 292294 149946 292874 149958
rect 328294 149946 328874 149958
rect 364294 149946 364874 149958
rect 400294 149946 400874 149958
rect 436294 149946 436874 149958
rect 472294 149946 472874 149958
rect 508294 149946 508874 149958
rect 544294 149946 544874 149958
rect 580294 149946 580874 149958
rect 587170 149946 587750 149958
rect -4746 149934 588670 149946
rect -4746 149698 -3654 149934
rect -3418 149698 4466 149934
rect 4702 149698 40466 149934
rect 40702 149698 76466 149934
rect 76702 149698 112466 149934
rect 112702 149698 148466 149934
rect 148702 149698 184466 149934
rect 184702 149698 220466 149934
rect 220702 149698 256466 149934
rect 256702 149698 292466 149934
rect 292702 149698 328466 149934
rect 328702 149698 364466 149934
rect 364702 149698 400466 149934
rect 400702 149698 436466 149934
rect 436702 149698 472466 149934
rect 472702 149698 508466 149934
rect 508702 149698 544466 149934
rect 544702 149698 580466 149934
rect 580702 149698 587342 149934
rect 587578 149698 588670 149934
rect -4746 149614 588670 149698
rect -4746 149378 -3654 149614
rect -3418 149378 4466 149614
rect 4702 149378 40466 149614
rect 40702 149378 76466 149614
rect 76702 149378 112466 149614
rect 112702 149378 148466 149614
rect 148702 149378 184466 149614
rect 184702 149378 220466 149614
rect 220702 149378 256466 149614
rect 256702 149378 292466 149614
rect 292702 149378 328466 149614
rect 328702 149378 364466 149614
rect 364702 149378 400466 149614
rect 400702 149378 436466 149614
rect 436702 149378 472466 149614
rect 472702 149378 508466 149614
rect 508702 149378 544466 149614
rect 544702 149378 580466 149614
rect 580702 149378 587342 149614
rect 587578 149378 588670 149614
rect -4746 149366 588670 149378
rect -3826 149354 -3246 149366
rect 4294 149354 4874 149366
rect 40294 149354 40874 149366
rect 76294 149354 76874 149366
rect 112294 149354 112874 149366
rect 148294 149354 148874 149366
rect 184294 149354 184874 149366
rect 220294 149354 220874 149366
rect 256294 149354 256874 149366
rect 292294 149354 292874 149366
rect 328294 149354 328874 149366
rect 364294 149354 364874 149366
rect 400294 149354 400874 149366
rect 436294 149354 436874 149366
rect 472294 149354 472874 149366
rect 508294 149354 508874 149366
rect 544294 149354 544874 149366
rect 580294 149354 580874 149366
rect 587170 149354 587750 149366
rect -1986 146466 -1406 146478
rect 814 146466 1394 146478
rect 36814 146466 37394 146478
rect 72814 146466 73394 146478
rect 108814 146466 109394 146478
rect 144814 146466 145394 146478
rect 180814 146466 181394 146478
rect 216814 146466 217394 146478
rect 252814 146466 253394 146478
rect 288814 146466 289394 146478
rect 324814 146466 325394 146478
rect 360814 146466 361394 146478
rect 396814 146466 397394 146478
rect 432814 146466 433394 146478
rect 468814 146466 469394 146478
rect 504814 146466 505394 146478
rect 540814 146466 541394 146478
rect 576814 146466 577394 146478
rect 585330 146466 585910 146478
rect -2906 146454 586830 146466
rect -2906 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586830 146454
rect -2906 146134 586830 146218
rect -2906 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586830 146134
rect -2906 145886 586830 145898
rect -1986 145874 -1406 145886
rect 814 145874 1394 145886
rect 36814 145874 37394 145886
rect 72814 145874 73394 145886
rect 108814 145874 109394 145886
rect 144814 145874 145394 145886
rect 180814 145874 181394 145886
rect 216814 145874 217394 145886
rect 252814 145874 253394 145886
rect 288814 145874 289394 145886
rect 324814 145874 325394 145886
rect 360814 145874 361394 145886
rect 396814 145874 397394 145886
rect 432814 145874 433394 145886
rect 468814 145874 469394 145886
rect 504814 145874 505394 145886
rect 540814 145874 541394 145886
rect 576814 145874 577394 145886
rect 585330 145874 585910 145886
rect -8426 138906 -7846 138918
rect 29254 138906 29834 138918
rect 65254 138906 65834 138918
rect 101254 138906 101834 138918
rect 137254 138906 137834 138918
rect 173254 138906 173834 138918
rect 209254 138906 209834 138918
rect 245254 138906 245834 138918
rect 281254 138906 281834 138918
rect 317254 138906 317834 138918
rect 353254 138906 353834 138918
rect 389254 138906 389834 138918
rect 425254 138906 425834 138918
rect 461254 138906 461834 138918
rect 497254 138906 497834 138918
rect 533254 138906 533834 138918
rect 569254 138906 569834 138918
rect 591770 138906 592350 138918
rect -8426 138894 592350 138906
rect -8426 138658 -8254 138894
rect -8018 138658 29426 138894
rect 29662 138658 65426 138894
rect 65662 138658 101426 138894
rect 101662 138658 137426 138894
rect 137662 138658 173426 138894
rect 173662 138658 209426 138894
rect 209662 138658 245426 138894
rect 245662 138658 281426 138894
rect 281662 138658 317426 138894
rect 317662 138658 353426 138894
rect 353662 138658 389426 138894
rect 389662 138658 425426 138894
rect 425662 138658 461426 138894
rect 461662 138658 497426 138894
rect 497662 138658 533426 138894
rect 533662 138658 569426 138894
rect 569662 138658 591942 138894
rect 592178 138658 592350 138894
rect -8426 138574 592350 138658
rect -8426 138338 -8254 138574
rect -8018 138338 29426 138574
rect 29662 138338 65426 138574
rect 65662 138338 101426 138574
rect 101662 138338 137426 138574
rect 137662 138338 173426 138574
rect 173662 138338 209426 138574
rect 209662 138338 245426 138574
rect 245662 138338 281426 138574
rect 281662 138338 317426 138574
rect 317662 138338 353426 138574
rect 353662 138338 389426 138574
rect 389662 138338 425426 138574
rect 425662 138338 461426 138574
rect 461662 138338 497426 138574
rect 497662 138338 533426 138574
rect 533662 138338 569426 138574
rect 569662 138338 591942 138574
rect 592178 138338 592350 138574
rect -8426 138326 592350 138338
rect -8426 138314 -7846 138326
rect 29254 138314 29834 138326
rect 65254 138314 65834 138326
rect 101254 138314 101834 138326
rect 137254 138314 137834 138326
rect 173254 138314 173834 138326
rect 209254 138314 209834 138326
rect 245254 138314 245834 138326
rect 281254 138314 281834 138326
rect 317254 138314 317834 138326
rect 353254 138314 353834 138326
rect 389254 138314 389834 138326
rect 425254 138314 425834 138326
rect 461254 138314 461834 138326
rect 497254 138314 497834 138326
rect 533254 138314 533834 138326
rect 569254 138314 569834 138326
rect 591770 138314 592350 138326
rect -6586 135426 -6006 135438
rect 25774 135426 26354 135438
rect 61774 135426 62354 135438
rect 97774 135426 98354 135438
rect 133774 135426 134354 135438
rect 169774 135426 170354 135438
rect 205774 135426 206354 135438
rect 241774 135426 242354 135438
rect 277774 135426 278354 135438
rect 313774 135426 314354 135438
rect 349774 135426 350354 135438
rect 385774 135426 386354 135438
rect 421774 135426 422354 135438
rect 457774 135426 458354 135438
rect 493774 135426 494354 135438
rect 529774 135426 530354 135438
rect 565774 135426 566354 135438
rect 589930 135426 590510 135438
rect -6586 135414 590510 135426
rect -6586 135178 -6414 135414
rect -6178 135178 25946 135414
rect 26182 135178 61946 135414
rect 62182 135178 97946 135414
rect 98182 135178 133946 135414
rect 134182 135178 169946 135414
rect 170182 135178 205946 135414
rect 206182 135178 241946 135414
rect 242182 135178 277946 135414
rect 278182 135178 313946 135414
rect 314182 135178 349946 135414
rect 350182 135178 385946 135414
rect 386182 135178 421946 135414
rect 422182 135178 457946 135414
rect 458182 135178 493946 135414
rect 494182 135178 529946 135414
rect 530182 135178 565946 135414
rect 566182 135178 590102 135414
rect 590338 135178 590510 135414
rect -6586 135094 590510 135178
rect -6586 134858 -6414 135094
rect -6178 134858 25946 135094
rect 26182 134858 61946 135094
rect 62182 134858 97946 135094
rect 98182 134858 133946 135094
rect 134182 134858 169946 135094
rect 170182 134858 205946 135094
rect 206182 134858 241946 135094
rect 242182 134858 277946 135094
rect 278182 134858 313946 135094
rect 314182 134858 349946 135094
rect 350182 134858 385946 135094
rect 386182 134858 421946 135094
rect 422182 134858 457946 135094
rect 458182 134858 493946 135094
rect 494182 134858 529946 135094
rect 530182 134858 565946 135094
rect 566182 134858 590102 135094
rect 590338 134858 590510 135094
rect -6586 134846 590510 134858
rect -6586 134834 -6006 134846
rect 25774 134834 26354 134846
rect 61774 134834 62354 134846
rect 97774 134834 98354 134846
rect 133774 134834 134354 134846
rect 169774 134834 170354 134846
rect 205774 134834 206354 134846
rect 241774 134834 242354 134846
rect 277774 134834 278354 134846
rect 313774 134834 314354 134846
rect 349774 134834 350354 134846
rect 385774 134834 386354 134846
rect 421774 134834 422354 134846
rect 457774 134834 458354 134846
rect 493774 134834 494354 134846
rect 529774 134834 530354 134846
rect 565774 134834 566354 134846
rect 589930 134834 590510 134846
rect -4746 131946 -4166 131958
rect 22294 131946 22874 131958
rect 58294 131946 58874 131958
rect 94294 131946 94874 131958
rect 130294 131946 130874 131958
rect 166294 131946 166874 131958
rect 202294 131946 202874 131958
rect 238294 131946 238874 131958
rect 274294 131946 274874 131958
rect 310294 131946 310874 131958
rect 346294 131946 346874 131958
rect 382294 131946 382874 131958
rect 418294 131946 418874 131958
rect 454294 131946 454874 131958
rect 490294 131946 490874 131958
rect 526294 131946 526874 131958
rect 562294 131946 562874 131958
rect 588090 131946 588670 131958
rect -4746 131934 588670 131946
rect -4746 131698 -4574 131934
rect -4338 131698 22466 131934
rect 22702 131698 58466 131934
rect 58702 131698 94466 131934
rect 94702 131698 130466 131934
rect 130702 131698 166466 131934
rect 166702 131698 202466 131934
rect 202702 131698 238466 131934
rect 238702 131698 274466 131934
rect 274702 131698 310466 131934
rect 310702 131698 346466 131934
rect 346702 131698 382466 131934
rect 382702 131698 418466 131934
rect 418702 131698 454466 131934
rect 454702 131698 490466 131934
rect 490702 131698 526466 131934
rect 526702 131698 562466 131934
rect 562702 131698 588262 131934
rect 588498 131698 588670 131934
rect -4746 131614 588670 131698
rect -4746 131378 -4574 131614
rect -4338 131378 22466 131614
rect 22702 131378 58466 131614
rect 58702 131378 94466 131614
rect 94702 131378 130466 131614
rect 130702 131378 166466 131614
rect 166702 131378 202466 131614
rect 202702 131378 238466 131614
rect 238702 131378 274466 131614
rect 274702 131378 310466 131614
rect 310702 131378 346466 131614
rect 346702 131378 382466 131614
rect 382702 131378 418466 131614
rect 418702 131378 454466 131614
rect 454702 131378 490466 131614
rect 490702 131378 526466 131614
rect 526702 131378 562466 131614
rect 562702 131378 588262 131614
rect 588498 131378 588670 131614
rect -4746 131366 588670 131378
rect -4746 131354 -4166 131366
rect 22294 131354 22874 131366
rect 58294 131354 58874 131366
rect 94294 131354 94874 131366
rect 130294 131354 130874 131366
rect 166294 131354 166874 131366
rect 202294 131354 202874 131366
rect 238294 131354 238874 131366
rect 274294 131354 274874 131366
rect 310294 131354 310874 131366
rect 346294 131354 346874 131366
rect 382294 131354 382874 131366
rect 418294 131354 418874 131366
rect 454294 131354 454874 131366
rect 490294 131354 490874 131366
rect 526294 131354 526874 131366
rect 562294 131354 562874 131366
rect 588090 131354 588670 131366
rect -2906 128466 -2326 128478
rect 18814 128466 19394 128478
rect 54814 128466 55394 128478
rect 90814 128466 91394 128478
rect 126814 128466 127394 128478
rect 162814 128466 163394 128478
rect 198814 128466 199394 128478
rect 234814 128466 235394 128478
rect 270814 128466 271394 128478
rect 306814 128466 307394 128478
rect 342814 128466 343394 128478
rect 378814 128466 379394 128478
rect 414814 128466 415394 128478
rect 450814 128466 451394 128478
rect 486814 128466 487394 128478
rect 522814 128466 523394 128478
rect 558814 128466 559394 128478
rect 586250 128466 586830 128478
rect -2906 128454 586830 128466
rect -2906 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586830 128454
rect -2906 128134 586830 128218
rect -2906 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586830 128134
rect -2906 127886 586830 127898
rect -2906 127874 -2326 127886
rect 18814 127874 19394 127886
rect 54814 127874 55394 127886
rect 90814 127874 91394 127886
rect 126814 127874 127394 127886
rect 162814 127874 163394 127886
rect 198814 127874 199394 127886
rect 234814 127874 235394 127886
rect 270814 127874 271394 127886
rect 306814 127874 307394 127886
rect 342814 127874 343394 127886
rect 378814 127874 379394 127886
rect 414814 127874 415394 127886
rect 450814 127874 451394 127886
rect 486814 127874 487394 127886
rect 522814 127874 523394 127886
rect 558814 127874 559394 127886
rect 586250 127874 586830 127886
rect -7506 120906 -6926 120918
rect 11254 120906 11834 120918
rect 47254 120906 47834 120918
rect 83254 120906 83834 120918
rect 119254 120906 119834 120918
rect 155254 120906 155834 120918
rect 191254 120906 191834 120918
rect 227254 120906 227834 120918
rect 263254 120906 263834 120918
rect 299254 120906 299834 120918
rect 335254 120906 335834 120918
rect 371254 120906 371834 120918
rect 407254 120906 407834 120918
rect 443254 120906 443834 120918
rect 479254 120906 479834 120918
rect 515254 120906 515834 120918
rect 551254 120906 551834 120918
rect 590850 120906 591430 120918
rect -8426 120894 592350 120906
rect -8426 120658 -7334 120894
rect -7098 120658 11426 120894
rect 11662 120658 47426 120894
rect 47662 120658 83426 120894
rect 83662 120658 119426 120894
rect 119662 120658 155426 120894
rect 155662 120658 191426 120894
rect 191662 120658 227426 120894
rect 227662 120658 263426 120894
rect 263662 120658 299426 120894
rect 299662 120658 335426 120894
rect 335662 120658 371426 120894
rect 371662 120658 407426 120894
rect 407662 120658 443426 120894
rect 443662 120658 479426 120894
rect 479662 120658 515426 120894
rect 515662 120658 551426 120894
rect 551662 120658 591022 120894
rect 591258 120658 592350 120894
rect -8426 120574 592350 120658
rect -8426 120338 -7334 120574
rect -7098 120338 11426 120574
rect 11662 120338 47426 120574
rect 47662 120338 83426 120574
rect 83662 120338 119426 120574
rect 119662 120338 155426 120574
rect 155662 120338 191426 120574
rect 191662 120338 227426 120574
rect 227662 120338 263426 120574
rect 263662 120338 299426 120574
rect 299662 120338 335426 120574
rect 335662 120338 371426 120574
rect 371662 120338 407426 120574
rect 407662 120338 443426 120574
rect 443662 120338 479426 120574
rect 479662 120338 515426 120574
rect 515662 120338 551426 120574
rect 551662 120338 591022 120574
rect 591258 120338 592350 120574
rect -8426 120326 592350 120338
rect -7506 120314 -6926 120326
rect 11254 120314 11834 120326
rect 47254 120314 47834 120326
rect 83254 120314 83834 120326
rect 119254 120314 119834 120326
rect 155254 120314 155834 120326
rect 191254 120314 191834 120326
rect 227254 120314 227834 120326
rect 263254 120314 263834 120326
rect 299254 120314 299834 120326
rect 335254 120314 335834 120326
rect 371254 120314 371834 120326
rect 407254 120314 407834 120326
rect 443254 120314 443834 120326
rect 479254 120314 479834 120326
rect 515254 120314 515834 120326
rect 551254 120314 551834 120326
rect 590850 120314 591430 120326
rect -5666 117426 -5086 117438
rect 7774 117426 8354 117438
rect 43774 117426 44354 117438
rect 79774 117426 80354 117438
rect 115774 117426 116354 117438
rect 151774 117426 152354 117438
rect 187774 117426 188354 117438
rect 223774 117426 224354 117438
rect 259774 117426 260354 117438
rect 295774 117426 296354 117438
rect 331774 117426 332354 117438
rect 367774 117426 368354 117438
rect 403774 117426 404354 117438
rect 439774 117426 440354 117438
rect 475774 117426 476354 117438
rect 511774 117426 512354 117438
rect 547774 117426 548354 117438
rect 589010 117426 589590 117438
rect -6586 117414 590510 117426
rect -6586 117178 -5494 117414
rect -5258 117178 7946 117414
rect 8182 117178 43946 117414
rect 44182 117178 79946 117414
rect 80182 117178 115946 117414
rect 116182 117178 151946 117414
rect 152182 117178 187946 117414
rect 188182 117178 223946 117414
rect 224182 117178 259946 117414
rect 260182 117178 295946 117414
rect 296182 117178 331946 117414
rect 332182 117178 367946 117414
rect 368182 117178 403946 117414
rect 404182 117178 439946 117414
rect 440182 117178 475946 117414
rect 476182 117178 511946 117414
rect 512182 117178 547946 117414
rect 548182 117178 589182 117414
rect 589418 117178 590510 117414
rect -6586 117094 590510 117178
rect -6586 116858 -5494 117094
rect -5258 116858 7946 117094
rect 8182 116858 43946 117094
rect 44182 116858 79946 117094
rect 80182 116858 115946 117094
rect 116182 116858 151946 117094
rect 152182 116858 187946 117094
rect 188182 116858 223946 117094
rect 224182 116858 259946 117094
rect 260182 116858 295946 117094
rect 296182 116858 331946 117094
rect 332182 116858 367946 117094
rect 368182 116858 403946 117094
rect 404182 116858 439946 117094
rect 440182 116858 475946 117094
rect 476182 116858 511946 117094
rect 512182 116858 547946 117094
rect 548182 116858 589182 117094
rect 589418 116858 590510 117094
rect -6586 116846 590510 116858
rect -5666 116834 -5086 116846
rect 7774 116834 8354 116846
rect 43774 116834 44354 116846
rect 79774 116834 80354 116846
rect 115774 116834 116354 116846
rect 151774 116834 152354 116846
rect 187774 116834 188354 116846
rect 223774 116834 224354 116846
rect 259774 116834 260354 116846
rect 295774 116834 296354 116846
rect 331774 116834 332354 116846
rect 367774 116834 368354 116846
rect 403774 116834 404354 116846
rect 439774 116834 440354 116846
rect 475774 116834 476354 116846
rect 511774 116834 512354 116846
rect 547774 116834 548354 116846
rect 589010 116834 589590 116846
rect -3826 113946 -3246 113958
rect 4294 113946 4874 113958
rect 40294 113946 40874 113958
rect 76294 113946 76874 113958
rect 112294 113946 112874 113958
rect 148294 113946 148874 113958
rect 184294 113946 184874 113958
rect 220294 113946 220874 113958
rect 256294 113946 256874 113958
rect 292294 113946 292874 113958
rect 328294 113946 328874 113958
rect 364294 113946 364874 113958
rect 400294 113946 400874 113958
rect 436294 113946 436874 113958
rect 472294 113946 472874 113958
rect 508294 113946 508874 113958
rect 544294 113946 544874 113958
rect 580294 113946 580874 113958
rect 587170 113946 587750 113958
rect -4746 113934 588670 113946
rect -4746 113698 -3654 113934
rect -3418 113698 4466 113934
rect 4702 113698 40466 113934
rect 40702 113698 76466 113934
rect 76702 113698 112466 113934
rect 112702 113698 148466 113934
rect 148702 113698 184466 113934
rect 184702 113698 220466 113934
rect 220702 113698 256466 113934
rect 256702 113698 292466 113934
rect 292702 113698 328466 113934
rect 328702 113698 364466 113934
rect 364702 113698 400466 113934
rect 400702 113698 436466 113934
rect 436702 113698 472466 113934
rect 472702 113698 508466 113934
rect 508702 113698 544466 113934
rect 544702 113698 580466 113934
rect 580702 113698 587342 113934
rect 587578 113698 588670 113934
rect -4746 113614 588670 113698
rect -4746 113378 -3654 113614
rect -3418 113378 4466 113614
rect 4702 113378 40466 113614
rect 40702 113378 76466 113614
rect 76702 113378 112466 113614
rect 112702 113378 148466 113614
rect 148702 113378 184466 113614
rect 184702 113378 220466 113614
rect 220702 113378 256466 113614
rect 256702 113378 292466 113614
rect 292702 113378 328466 113614
rect 328702 113378 364466 113614
rect 364702 113378 400466 113614
rect 400702 113378 436466 113614
rect 436702 113378 472466 113614
rect 472702 113378 508466 113614
rect 508702 113378 544466 113614
rect 544702 113378 580466 113614
rect 580702 113378 587342 113614
rect 587578 113378 588670 113614
rect -4746 113366 588670 113378
rect -3826 113354 -3246 113366
rect 4294 113354 4874 113366
rect 40294 113354 40874 113366
rect 76294 113354 76874 113366
rect 112294 113354 112874 113366
rect 148294 113354 148874 113366
rect 184294 113354 184874 113366
rect 220294 113354 220874 113366
rect 256294 113354 256874 113366
rect 292294 113354 292874 113366
rect 328294 113354 328874 113366
rect 364294 113354 364874 113366
rect 400294 113354 400874 113366
rect 436294 113354 436874 113366
rect 472294 113354 472874 113366
rect 508294 113354 508874 113366
rect 544294 113354 544874 113366
rect 580294 113354 580874 113366
rect 587170 113354 587750 113366
rect -1986 110466 -1406 110478
rect 814 110466 1394 110478
rect 36814 110466 37394 110478
rect 72814 110466 73394 110478
rect 108814 110466 109394 110478
rect 144814 110466 145394 110478
rect 180814 110466 181394 110478
rect 216814 110466 217394 110478
rect 252814 110466 253394 110478
rect 288814 110466 289394 110478
rect 324814 110466 325394 110478
rect 360814 110466 361394 110478
rect 396814 110466 397394 110478
rect 432814 110466 433394 110478
rect 468814 110466 469394 110478
rect 504814 110466 505394 110478
rect 540814 110466 541394 110478
rect 576814 110466 577394 110478
rect 585330 110466 585910 110478
rect -2906 110454 586830 110466
rect -2906 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586830 110454
rect -2906 110134 586830 110218
rect -2906 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586830 110134
rect -2906 109886 586830 109898
rect -1986 109874 -1406 109886
rect 814 109874 1394 109886
rect 36814 109874 37394 109886
rect 72814 109874 73394 109886
rect 108814 109874 109394 109886
rect 144814 109874 145394 109886
rect 180814 109874 181394 109886
rect 216814 109874 217394 109886
rect 252814 109874 253394 109886
rect 288814 109874 289394 109886
rect 324814 109874 325394 109886
rect 360814 109874 361394 109886
rect 396814 109874 397394 109886
rect 432814 109874 433394 109886
rect 468814 109874 469394 109886
rect 504814 109874 505394 109886
rect 540814 109874 541394 109886
rect 576814 109874 577394 109886
rect 585330 109874 585910 109886
rect -8426 102906 -7846 102918
rect 29254 102906 29834 102918
rect 65254 102906 65834 102918
rect 101254 102906 101834 102918
rect 137254 102906 137834 102918
rect 173254 102906 173834 102918
rect 209254 102906 209834 102918
rect 245254 102906 245834 102918
rect 281254 102906 281834 102918
rect 317254 102906 317834 102918
rect 353254 102906 353834 102918
rect 389254 102906 389834 102918
rect 425254 102906 425834 102918
rect 461254 102906 461834 102918
rect 497254 102906 497834 102918
rect 533254 102906 533834 102918
rect 569254 102906 569834 102918
rect 591770 102906 592350 102918
rect -8426 102894 592350 102906
rect -8426 102658 -8254 102894
rect -8018 102658 29426 102894
rect 29662 102658 65426 102894
rect 65662 102658 101426 102894
rect 101662 102658 137426 102894
rect 137662 102658 173426 102894
rect 173662 102658 209426 102894
rect 209662 102658 245426 102894
rect 245662 102658 281426 102894
rect 281662 102658 317426 102894
rect 317662 102658 353426 102894
rect 353662 102658 389426 102894
rect 389662 102658 425426 102894
rect 425662 102658 461426 102894
rect 461662 102658 497426 102894
rect 497662 102658 533426 102894
rect 533662 102658 569426 102894
rect 569662 102658 591942 102894
rect 592178 102658 592350 102894
rect -8426 102574 592350 102658
rect -8426 102338 -8254 102574
rect -8018 102338 29426 102574
rect 29662 102338 65426 102574
rect 65662 102338 101426 102574
rect 101662 102338 137426 102574
rect 137662 102338 173426 102574
rect 173662 102338 209426 102574
rect 209662 102338 245426 102574
rect 245662 102338 281426 102574
rect 281662 102338 317426 102574
rect 317662 102338 353426 102574
rect 353662 102338 389426 102574
rect 389662 102338 425426 102574
rect 425662 102338 461426 102574
rect 461662 102338 497426 102574
rect 497662 102338 533426 102574
rect 533662 102338 569426 102574
rect 569662 102338 591942 102574
rect 592178 102338 592350 102574
rect -8426 102326 592350 102338
rect -8426 102314 -7846 102326
rect 29254 102314 29834 102326
rect 65254 102314 65834 102326
rect 101254 102314 101834 102326
rect 137254 102314 137834 102326
rect 173254 102314 173834 102326
rect 209254 102314 209834 102326
rect 245254 102314 245834 102326
rect 281254 102314 281834 102326
rect 317254 102314 317834 102326
rect 353254 102314 353834 102326
rect 389254 102314 389834 102326
rect 425254 102314 425834 102326
rect 461254 102314 461834 102326
rect 497254 102314 497834 102326
rect 533254 102314 533834 102326
rect 569254 102314 569834 102326
rect 591770 102314 592350 102326
rect -6586 99426 -6006 99438
rect 25774 99426 26354 99438
rect 61774 99426 62354 99438
rect 97774 99426 98354 99438
rect 133774 99426 134354 99438
rect 169774 99426 170354 99438
rect 205774 99426 206354 99438
rect 241774 99426 242354 99438
rect 277774 99426 278354 99438
rect 313774 99426 314354 99438
rect 349774 99426 350354 99438
rect 385774 99426 386354 99438
rect 421774 99426 422354 99438
rect 457774 99426 458354 99438
rect 493774 99426 494354 99438
rect 529774 99426 530354 99438
rect 565774 99426 566354 99438
rect 589930 99426 590510 99438
rect -6586 99414 590510 99426
rect -6586 99178 -6414 99414
rect -6178 99178 25946 99414
rect 26182 99178 61946 99414
rect 62182 99178 97946 99414
rect 98182 99178 133946 99414
rect 134182 99178 169946 99414
rect 170182 99178 205946 99414
rect 206182 99178 241946 99414
rect 242182 99178 277946 99414
rect 278182 99178 313946 99414
rect 314182 99178 349946 99414
rect 350182 99178 385946 99414
rect 386182 99178 421946 99414
rect 422182 99178 457946 99414
rect 458182 99178 493946 99414
rect 494182 99178 529946 99414
rect 530182 99178 565946 99414
rect 566182 99178 590102 99414
rect 590338 99178 590510 99414
rect -6586 99094 590510 99178
rect -6586 98858 -6414 99094
rect -6178 98858 25946 99094
rect 26182 98858 61946 99094
rect 62182 98858 97946 99094
rect 98182 98858 133946 99094
rect 134182 98858 169946 99094
rect 170182 98858 205946 99094
rect 206182 98858 241946 99094
rect 242182 98858 277946 99094
rect 278182 98858 313946 99094
rect 314182 98858 349946 99094
rect 350182 98858 385946 99094
rect 386182 98858 421946 99094
rect 422182 98858 457946 99094
rect 458182 98858 493946 99094
rect 494182 98858 529946 99094
rect 530182 98858 565946 99094
rect 566182 98858 590102 99094
rect 590338 98858 590510 99094
rect -6586 98846 590510 98858
rect -6586 98834 -6006 98846
rect 25774 98834 26354 98846
rect 61774 98834 62354 98846
rect 97774 98834 98354 98846
rect 133774 98834 134354 98846
rect 169774 98834 170354 98846
rect 205774 98834 206354 98846
rect 241774 98834 242354 98846
rect 277774 98834 278354 98846
rect 313774 98834 314354 98846
rect 349774 98834 350354 98846
rect 385774 98834 386354 98846
rect 421774 98834 422354 98846
rect 457774 98834 458354 98846
rect 493774 98834 494354 98846
rect 529774 98834 530354 98846
rect 565774 98834 566354 98846
rect 589930 98834 590510 98846
rect -4746 95946 -4166 95958
rect 22294 95946 22874 95958
rect 58294 95946 58874 95958
rect 94294 95946 94874 95958
rect 130294 95946 130874 95958
rect 166294 95946 166874 95958
rect 202294 95946 202874 95958
rect 238294 95946 238874 95958
rect 274294 95946 274874 95958
rect 310294 95946 310874 95958
rect 346294 95946 346874 95958
rect 382294 95946 382874 95958
rect 418294 95946 418874 95958
rect 454294 95946 454874 95958
rect 490294 95946 490874 95958
rect 526294 95946 526874 95958
rect 562294 95946 562874 95958
rect 588090 95946 588670 95958
rect -4746 95934 588670 95946
rect -4746 95698 -4574 95934
rect -4338 95698 22466 95934
rect 22702 95698 58466 95934
rect 58702 95698 94466 95934
rect 94702 95698 130466 95934
rect 130702 95698 166466 95934
rect 166702 95698 202466 95934
rect 202702 95698 238466 95934
rect 238702 95698 274466 95934
rect 274702 95698 310466 95934
rect 310702 95698 346466 95934
rect 346702 95698 382466 95934
rect 382702 95698 418466 95934
rect 418702 95698 454466 95934
rect 454702 95698 490466 95934
rect 490702 95698 526466 95934
rect 526702 95698 562466 95934
rect 562702 95698 588262 95934
rect 588498 95698 588670 95934
rect -4746 95614 588670 95698
rect -4746 95378 -4574 95614
rect -4338 95378 22466 95614
rect 22702 95378 58466 95614
rect 58702 95378 94466 95614
rect 94702 95378 130466 95614
rect 130702 95378 166466 95614
rect 166702 95378 202466 95614
rect 202702 95378 238466 95614
rect 238702 95378 274466 95614
rect 274702 95378 310466 95614
rect 310702 95378 346466 95614
rect 346702 95378 382466 95614
rect 382702 95378 418466 95614
rect 418702 95378 454466 95614
rect 454702 95378 490466 95614
rect 490702 95378 526466 95614
rect 526702 95378 562466 95614
rect 562702 95378 588262 95614
rect 588498 95378 588670 95614
rect -4746 95366 588670 95378
rect -4746 95354 -4166 95366
rect 22294 95354 22874 95366
rect 58294 95354 58874 95366
rect 94294 95354 94874 95366
rect 130294 95354 130874 95366
rect 166294 95354 166874 95366
rect 202294 95354 202874 95366
rect 238294 95354 238874 95366
rect 274294 95354 274874 95366
rect 310294 95354 310874 95366
rect 346294 95354 346874 95366
rect 382294 95354 382874 95366
rect 418294 95354 418874 95366
rect 454294 95354 454874 95366
rect 490294 95354 490874 95366
rect 526294 95354 526874 95366
rect 562294 95354 562874 95366
rect 588090 95354 588670 95366
rect -2906 92466 -2326 92478
rect 18814 92466 19394 92478
rect 54814 92466 55394 92478
rect 90814 92466 91394 92478
rect 126814 92466 127394 92478
rect 162814 92466 163394 92478
rect 198814 92466 199394 92478
rect 234814 92466 235394 92478
rect 270814 92466 271394 92478
rect 306814 92466 307394 92478
rect 342814 92466 343394 92478
rect 378814 92466 379394 92478
rect 414814 92466 415394 92478
rect 450814 92466 451394 92478
rect 486814 92466 487394 92478
rect 522814 92466 523394 92478
rect 558814 92466 559394 92478
rect 586250 92466 586830 92478
rect -2906 92454 586830 92466
rect -2906 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586830 92454
rect -2906 92134 586830 92218
rect -2906 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586830 92134
rect -2906 91886 586830 91898
rect -2906 91874 -2326 91886
rect 18814 91874 19394 91886
rect 54814 91874 55394 91886
rect 90814 91874 91394 91886
rect 126814 91874 127394 91886
rect 162814 91874 163394 91886
rect 198814 91874 199394 91886
rect 234814 91874 235394 91886
rect 270814 91874 271394 91886
rect 306814 91874 307394 91886
rect 342814 91874 343394 91886
rect 378814 91874 379394 91886
rect 414814 91874 415394 91886
rect 450814 91874 451394 91886
rect 486814 91874 487394 91886
rect 522814 91874 523394 91886
rect 558814 91874 559394 91886
rect 586250 91874 586830 91886
rect -7506 84906 -6926 84918
rect 11254 84906 11834 84918
rect 47254 84906 47834 84918
rect 83254 84906 83834 84918
rect 119254 84906 119834 84918
rect 155254 84906 155834 84918
rect 191254 84906 191834 84918
rect 227254 84906 227834 84918
rect 263254 84906 263834 84918
rect 299254 84906 299834 84918
rect 335254 84906 335834 84918
rect 371254 84906 371834 84918
rect 407254 84906 407834 84918
rect 443254 84906 443834 84918
rect 479254 84906 479834 84918
rect 515254 84906 515834 84918
rect 551254 84906 551834 84918
rect 590850 84906 591430 84918
rect -8426 84894 592350 84906
rect -8426 84658 -7334 84894
rect -7098 84658 11426 84894
rect 11662 84658 47426 84894
rect 47662 84658 83426 84894
rect 83662 84658 119426 84894
rect 119662 84658 155426 84894
rect 155662 84658 191426 84894
rect 191662 84658 227426 84894
rect 227662 84658 263426 84894
rect 263662 84658 299426 84894
rect 299662 84658 335426 84894
rect 335662 84658 371426 84894
rect 371662 84658 407426 84894
rect 407662 84658 443426 84894
rect 443662 84658 479426 84894
rect 479662 84658 515426 84894
rect 515662 84658 551426 84894
rect 551662 84658 591022 84894
rect 591258 84658 592350 84894
rect -8426 84574 592350 84658
rect -8426 84338 -7334 84574
rect -7098 84338 11426 84574
rect 11662 84338 47426 84574
rect 47662 84338 83426 84574
rect 83662 84338 119426 84574
rect 119662 84338 155426 84574
rect 155662 84338 191426 84574
rect 191662 84338 227426 84574
rect 227662 84338 263426 84574
rect 263662 84338 299426 84574
rect 299662 84338 335426 84574
rect 335662 84338 371426 84574
rect 371662 84338 407426 84574
rect 407662 84338 443426 84574
rect 443662 84338 479426 84574
rect 479662 84338 515426 84574
rect 515662 84338 551426 84574
rect 551662 84338 591022 84574
rect 591258 84338 592350 84574
rect -8426 84326 592350 84338
rect -7506 84314 -6926 84326
rect 11254 84314 11834 84326
rect 47254 84314 47834 84326
rect 83254 84314 83834 84326
rect 119254 84314 119834 84326
rect 155254 84314 155834 84326
rect 191254 84314 191834 84326
rect 227254 84314 227834 84326
rect 263254 84314 263834 84326
rect 299254 84314 299834 84326
rect 335254 84314 335834 84326
rect 371254 84314 371834 84326
rect 407254 84314 407834 84326
rect 443254 84314 443834 84326
rect 479254 84314 479834 84326
rect 515254 84314 515834 84326
rect 551254 84314 551834 84326
rect 590850 84314 591430 84326
rect -5666 81426 -5086 81438
rect 7774 81426 8354 81438
rect 43774 81426 44354 81438
rect 79774 81426 80354 81438
rect 115774 81426 116354 81438
rect 151774 81426 152354 81438
rect 187774 81426 188354 81438
rect 223774 81426 224354 81438
rect 259774 81426 260354 81438
rect 295774 81426 296354 81438
rect 331774 81426 332354 81438
rect 367774 81426 368354 81438
rect 403774 81426 404354 81438
rect 439774 81426 440354 81438
rect 475774 81426 476354 81438
rect 511774 81426 512354 81438
rect 547774 81426 548354 81438
rect 589010 81426 589590 81438
rect -6586 81414 590510 81426
rect -6586 81178 -5494 81414
rect -5258 81178 7946 81414
rect 8182 81178 43946 81414
rect 44182 81178 79946 81414
rect 80182 81178 115946 81414
rect 116182 81178 151946 81414
rect 152182 81178 187946 81414
rect 188182 81178 223946 81414
rect 224182 81178 259946 81414
rect 260182 81178 295946 81414
rect 296182 81178 331946 81414
rect 332182 81178 367946 81414
rect 368182 81178 403946 81414
rect 404182 81178 439946 81414
rect 440182 81178 475946 81414
rect 476182 81178 511946 81414
rect 512182 81178 547946 81414
rect 548182 81178 589182 81414
rect 589418 81178 590510 81414
rect -6586 81094 590510 81178
rect -6586 80858 -5494 81094
rect -5258 80858 7946 81094
rect 8182 80858 43946 81094
rect 44182 80858 79946 81094
rect 80182 80858 115946 81094
rect 116182 80858 151946 81094
rect 152182 80858 187946 81094
rect 188182 80858 223946 81094
rect 224182 80858 259946 81094
rect 260182 80858 295946 81094
rect 296182 80858 331946 81094
rect 332182 80858 367946 81094
rect 368182 80858 403946 81094
rect 404182 80858 439946 81094
rect 440182 80858 475946 81094
rect 476182 80858 511946 81094
rect 512182 80858 547946 81094
rect 548182 80858 589182 81094
rect 589418 80858 590510 81094
rect -6586 80846 590510 80858
rect -5666 80834 -5086 80846
rect 7774 80834 8354 80846
rect 43774 80834 44354 80846
rect 79774 80834 80354 80846
rect 115774 80834 116354 80846
rect 151774 80834 152354 80846
rect 187774 80834 188354 80846
rect 223774 80834 224354 80846
rect 259774 80834 260354 80846
rect 295774 80834 296354 80846
rect 331774 80834 332354 80846
rect 367774 80834 368354 80846
rect 403774 80834 404354 80846
rect 439774 80834 440354 80846
rect 475774 80834 476354 80846
rect 511774 80834 512354 80846
rect 547774 80834 548354 80846
rect 589010 80834 589590 80846
rect -3826 77946 -3246 77958
rect 4294 77946 4874 77958
rect 40294 77946 40874 77958
rect 76294 77946 76874 77958
rect 112294 77946 112874 77958
rect 148294 77946 148874 77958
rect 184294 77946 184874 77958
rect 220294 77946 220874 77958
rect 256294 77946 256874 77958
rect 292294 77946 292874 77958
rect 328294 77946 328874 77958
rect 364294 77946 364874 77958
rect 400294 77946 400874 77958
rect 436294 77946 436874 77958
rect 472294 77946 472874 77958
rect 508294 77946 508874 77958
rect 544294 77946 544874 77958
rect 580294 77946 580874 77958
rect 587170 77946 587750 77958
rect -4746 77934 588670 77946
rect -4746 77698 -3654 77934
rect -3418 77698 4466 77934
rect 4702 77698 40466 77934
rect 40702 77698 76466 77934
rect 76702 77698 112466 77934
rect 112702 77698 148466 77934
rect 148702 77698 184466 77934
rect 184702 77698 220466 77934
rect 220702 77698 256466 77934
rect 256702 77698 292466 77934
rect 292702 77698 328466 77934
rect 328702 77698 364466 77934
rect 364702 77698 400466 77934
rect 400702 77698 436466 77934
rect 436702 77698 472466 77934
rect 472702 77698 508466 77934
rect 508702 77698 544466 77934
rect 544702 77698 580466 77934
rect 580702 77698 587342 77934
rect 587578 77698 588670 77934
rect -4746 77614 588670 77698
rect -4746 77378 -3654 77614
rect -3418 77378 4466 77614
rect 4702 77378 40466 77614
rect 40702 77378 76466 77614
rect 76702 77378 112466 77614
rect 112702 77378 148466 77614
rect 148702 77378 184466 77614
rect 184702 77378 220466 77614
rect 220702 77378 256466 77614
rect 256702 77378 292466 77614
rect 292702 77378 328466 77614
rect 328702 77378 364466 77614
rect 364702 77378 400466 77614
rect 400702 77378 436466 77614
rect 436702 77378 472466 77614
rect 472702 77378 508466 77614
rect 508702 77378 544466 77614
rect 544702 77378 580466 77614
rect 580702 77378 587342 77614
rect 587578 77378 588670 77614
rect -4746 77366 588670 77378
rect -3826 77354 -3246 77366
rect 4294 77354 4874 77366
rect 40294 77354 40874 77366
rect 76294 77354 76874 77366
rect 112294 77354 112874 77366
rect 148294 77354 148874 77366
rect 184294 77354 184874 77366
rect 220294 77354 220874 77366
rect 256294 77354 256874 77366
rect 292294 77354 292874 77366
rect 328294 77354 328874 77366
rect 364294 77354 364874 77366
rect 400294 77354 400874 77366
rect 436294 77354 436874 77366
rect 472294 77354 472874 77366
rect 508294 77354 508874 77366
rect 544294 77354 544874 77366
rect 580294 77354 580874 77366
rect 587170 77354 587750 77366
rect -1986 74466 -1406 74478
rect 814 74466 1394 74478
rect 36814 74466 37394 74478
rect 72814 74466 73394 74478
rect 108814 74466 109394 74478
rect 144814 74466 145394 74478
rect 180814 74466 181394 74478
rect 216814 74466 217394 74478
rect 252814 74466 253394 74478
rect 288814 74466 289394 74478
rect 324814 74466 325394 74478
rect 360814 74466 361394 74478
rect 396814 74466 397394 74478
rect 432814 74466 433394 74478
rect 468814 74466 469394 74478
rect 504814 74466 505394 74478
rect 540814 74466 541394 74478
rect 576814 74466 577394 74478
rect 585330 74466 585910 74478
rect -2906 74454 586830 74466
rect -2906 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586830 74454
rect -2906 74134 586830 74218
rect -2906 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586830 74134
rect -2906 73886 586830 73898
rect -1986 73874 -1406 73886
rect 814 73874 1394 73886
rect 36814 73874 37394 73886
rect 72814 73874 73394 73886
rect 108814 73874 109394 73886
rect 144814 73874 145394 73886
rect 180814 73874 181394 73886
rect 216814 73874 217394 73886
rect 252814 73874 253394 73886
rect 288814 73874 289394 73886
rect 324814 73874 325394 73886
rect 360814 73874 361394 73886
rect 396814 73874 397394 73886
rect 432814 73874 433394 73886
rect 468814 73874 469394 73886
rect 504814 73874 505394 73886
rect 540814 73874 541394 73886
rect 576814 73874 577394 73886
rect 585330 73874 585910 73886
rect -8426 66906 -7846 66918
rect 29254 66906 29834 66918
rect 65254 66906 65834 66918
rect 101254 66906 101834 66918
rect 137254 66906 137834 66918
rect 173254 66906 173834 66918
rect 209254 66906 209834 66918
rect 245254 66906 245834 66918
rect 281254 66906 281834 66918
rect 317254 66906 317834 66918
rect 353254 66906 353834 66918
rect 389254 66906 389834 66918
rect 425254 66906 425834 66918
rect 461254 66906 461834 66918
rect 497254 66906 497834 66918
rect 533254 66906 533834 66918
rect 569254 66906 569834 66918
rect 591770 66906 592350 66918
rect -8426 66894 592350 66906
rect -8426 66658 -8254 66894
rect -8018 66658 29426 66894
rect 29662 66658 65426 66894
rect 65662 66658 101426 66894
rect 101662 66658 137426 66894
rect 137662 66658 173426 66894
rect 173662 66658 209426 66894
rect 209662 66658 245426 66894
rect 245662 66658 281426 66894
rect 281662 66658 317426 66894
rect 317662 66658 353426 66894
rect 353662 66658 389426 66894
rect 389662 66658 425426 66894
rect 425662 66658 461426 66894
rect 461662 66658 497426 66894
rect 497662 66658 533426 66894
rect 533662 66658 569426 66894
rect 569662 66658 591942 66894
rect 592178 66658 592350 66894
rect -8426 66574 592350 66658
rect -8426 66338 -8254 66574
rect -8018 66338 29426 66574
rect 29662 66338 65426 66574
rect 65662 66338 101426 66574
rect 101662 66338 137426 66574
rect 137662 66338 173426 66574
rect 173662 66338 209426 66574
rect 209662 66338 245426 66574
rect 245662 66338 281426 66574
rect 281662 66338 317426 66574
rect 317662 66338 353426 66574
rect 353662 66338 389426 66574
rect 389662 66338 425426 66574
rect 425662 66338 461426 66574
rect 461662 66338 497426 66574
rect 497662 66338 533426 66574
rect 533662 66338 569426 66574
rect 569662 66338 591942 66574
rect 592178 66338 592350 66574
rect -8426 66326 592350 66338
rect -8426 66314 -7846 66326
rect 29254 66314 29834 66326
rect 65254 66314 65834 66326
rect 101254 66314 101834 66326
rect 137254 66314 137834 66326
rect 173254 66314 173834 66326
rect 209254 66314 209834 66326
rect 245254 66314 245834 66326
rect 281254 66314 281834 66326
rect 317254 66314 317834 66326
rect 353254 66314 353834 66326
rect 389254 66314 389834 66326
rect 425254 66314 425834 66326
rect 461254 66314 461834 66326
rect 497254 66314 497834 66326
rect 533254 66314 533834 66326
rect 569254 66314 569834 66326
rect 591770 66314 592350 66326
rect -6586 63426 -6006 63438
rect 25774 63426 26354 63438
rect 61774 63426 62354 63438
rect 97774 63426 98354 63438
rect 133774 63426 134354 63438
rect 169774 63426 170354 63438
rect 205774 63426 206354 63438
rect 241774 63426 242354 63438
rect 277774 63426 278354 63438
rect 313774 63426 314354 63438
rect 349774 63426 350354 63438
rect 385774 63426 386354 63438
rect 421774 63426 422354 63438
rect 457774 63426 458354 63438
rect 493774 63426 494354 63438
rect 529774 63426 530354 63438
rect 565774 63426 566354 63438
rect 589930 63426 590510 63438
rect -6586 63414 590510 63426
rect -6586 63178 -6414 63414
rect -6178 63178 25946 63414
rect 26182 63178 61946 63414
rect 62182 63178 97946 63414
rect 98182 63178 133946 63414
rect 134182 63178 169946 63414
rect 170182 63178 205946 63414
rect 206182 63178 241946 63414
rect 242182 63178 277946 63414
rect 278182 63178 313946 63414
rect 314182 63178 349946 63414
rect 350182 63178 385946 63414
rect 386182 63178 421946 63414
rect 422182 63178 457946 63414
rect 458182 63178 493946 63414
rect 494182 63178 529946 63414
rect 530182 63178 565946 63414
rect 566182 63178 590102 63414
rect 590338 63178 590510 63414
rect -6586 63094 590510 63178
rect -6586 62858 -6414 63094
rect -6178 62858 25946 63094
rect 26182 62858 61946 63094
rect 62182 62858 97946 63094
rect 98182 62858 133946 63094
rect 134182 62858 169946 63094
rect 170182 62858 205946 63094
rect 206182 62858 241946 63094
rect 242182 62858 277946 63094
rect 278182 62858 313946 63094
rect 314182 62858 349946 63094
rect 350182 62858 385946 63094
rect 386182 62858 421946 63094
rect 422182 62858 457946 63094
rect 458182 62858 493946 63094
rect 494182 62858 529946 63094
rect 530182 62858 565946 63094
rect 566182 62858 590102 63094
rect 590338 62858 590510 63094
rect -6586 62846 590510 62858
rect -6586 62834 -6006 62846
rect 25774 62834 26354 62846
rect 61774 62834 62354 62846
rect 97774 62834 98354 62846
rect 133774 62834 134354 62846
rect 169774 62834 170354 62846
rect 205774 62834 206354 62846
rect 241774 62834 242354 62846
rect 277774 62834 278354 62846
rect 313774 62834 314354 62846
rect 349774 62834 350354 62846
rect 385774 62834 386354 62846
rect 421774 62834 422354 62846
rect 457774 62834 458354 62846
rect 493774 62834 494354 62846
rect 529774 62834 530354 62846
rect 565774 62834 566354 62846
rect 589930 62834 590510 62846
rect -4746 59946 -4166 59958
rect 22294 59946 22874 59958
rect 58294 59946 58874 59958
rect 94294 59946 94874 59958
rect 130294 59946 130874 59958
rect 166294 59946 166874 59958
rect 202294 59946 202874 59958
rect 238294 59946 238874 59958
rect 274294 59946 274874 59958
rect 310294 59946 310874 59958
rect 346294 59946 346874 59958
rect 382294 59946 382874 59958
rect 418294 59946 418874 59958
rect 454294 59946 454874 59958
rect 490294 59946 490874 59958
rect 526294 59946 526874 59958
rect 562294 59946 562874 59958
rect 588090 59946 588670 59958
rect -4746 59934 588670 59946
rect -4746 59698 -4574 59934
rect -4338 59698 22466 59934
rect 22702 59698 58466 59934
rect 58702 59698 94466 59934
rect 94702 59698 130466 59934
rect 130702 59698 166466 59934
rect 166702 59698 202466 59934
rect 202702 59698 238466 59934
rect 238702 59698 274466 59934
rect 274702 59698 310466 59934
rect 310702 59698 346466 59934
rect 346702 59698 382466 59934
rect 382702 59698 418466 59934
rect 418702 59698 454466 59934
rect 454702 59698 490466 59934
rect 490702 59698 526466 59934
rect 526702 59698 562466 59934
rect 562702 59698 588262 59934
rect 588498 59698 588670 59934
rect -4746 59614 588670 59698
rect -4746 59378 -4574 59614
rect -4338 59378 22466 59614
rect 22702 59378 58466 59614
rect 58702 59378 94466 59614
rect 94702 59378 130466 59614
rect 130702 59378 166466 59614
rect 166702 59378 202466 59614
rect 202702 59378 238466 59614
rect 238702 59378 274466 59614
rect 274702 59378 310466 59614
rect 310702 59378 346466 59614
rect 346702 59378 382466 59614
rect 382702 59378 418466 59614
rect 418702 59378 454466 59614
rect 454702 59378 490466 59614
rect 490702 59378 526466 59614
rect 526702 59378 562466 59614
rect 562702 59378 588262 59614
rect 588498 59378 588670 59614
rect -4746 59366 588670 59378
rect -4746 59354 -4166 59366
rect 22294 59354 22874 59366
rect 58294 59354 58874 59366
rect 94294 59354 94874 59366
rect 130294 59354 130874 59366
rect 166294 59354 166874 59366
rect 202294 59354 202874 59366
rect 238294 59354 238874 59366
rect 274294 59354 274874 59366
rect 310294 59354 310874 59366
rect 346294 59354 346874 59366
rect 382294 59354 382874 59366
rect 418294 59354 418874 59366
rect 454294 59354 454874 59366
rect 490294 59354 490874 59366
rect 526294 59354 526874 59366
rect 562294 59354 562874 59366
rect 588090 59354 588670 59366
rect -2906 56466 -2326 56478
rect 18814 56466 19394 56478
rect 54814 56466 55394 56478
rect 90814 56466 91394 56478
rect 126814 56466 127394 56478
rect 162814 56466 163394 56478
rect 198814 56466 199394 56478
rect 234814 56466 235394 56478
rect 270814 56466 271394 56478
rect 306814 56466 307394 56478
rect 342814 56466 343394 56478
rect 378814 56466 379394 56478
rect 414814 56466 415394 56478
rect 450814 56466 451394 56478
rect 486814 56466 487394 56478
rect 522814 56466 523394 56478
rect 558814 56466 559394 56478
rect 586250 56466 586830 56478
rect -2906 56454 586830 56466
rect -2906 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586830 56454
rect -2906 56134 586830 56218
rect -2906 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586830 56134
rect -2906 55886 586830 55898
rect -2906 55874 -2326 55886
rect 18814 55874 19394 55886
rect 54814 55874 55394 55886
rect 90814 55874 91394 55886
rect 126814 55874 127394 55886
rect 162814 55874 163394 55886
rect 198814 55874 199394 55886
rect 234814 55874 235394 55886
rect 270814 55874 271394 55886
rect 306814 55874 307394 55886
rect 342814 55874 343394 55886
rect 378814 55874 379394 55886
rect 414814 55874 415394 55886
rect 450814 55874 451394 55886
rect 486814 55874 487394 55886
rect 522814 55874 523394 55886
rect 558814 55874 559394 55886
rect 586250 55874 586830 55886
rect -7506 48906 -6926 48918
rect 11254 48906 11834 48918
rect 47254 48906 47834 48918
rect 83254 48906 83834 48918
rect 119254 48906 119834 48918
rect 155254 48906 155834 48918
rect 191254 48906 191834 48918
rect 227254 48906 227834 48918
rect 263254 48906 263834 48918
rect 299254 48906 299834 48918
rect 335254 48906 335834 48918
rect 371254 48906 371834 48918
rect 407254 48906 407834 48918
rect 443254 48906 443834 48918
rect 479254 48906 479834 48918
rect 515254 48906 515834 48918
rect 551254 48906 551834 48918
rect 590850 48906 591430 48918
rect -8426 48894 592350 48906
rect -8426 48658 -7334 48894
rect -7098 48658 11426 48894
rect 11662 48658 47426 48894
rect 47662 48658 83426 48894
rect 83662 48658 119426 48894
rect 119662 48658 155426 48894
rect 155662 48658 191426 48894
rect 191662 48658 227426 48894
rect 227662 48658 263426 48894
rect 263662 48658 299426 48894
rect 299662 48658 335426 48894
rect 335662 48658 371426 48894
rect 371662 48658 407426 48894
rect 407662 48658 443426 48894
rect 443662 48658 479426 48894
rect 479662 48658 515426 48894
rect 515662 48658 551426 48894
rect 551662 48658 591022 48894
rect 591258 48658 592350 48894
rect -8426 48574 592350 48658
rect -8426 48338 -7334 48574
rect -7098 48338 11426 48574
rect 11662 48338 47426 48574
rect 47662 48338 83426 48574
rect 83662 48338 119426 48574
rect 119662 48338 155426 48574
rect 155662 48338 191426 48574
rect 191662 48338 227426 48574
rect 227662 48338 263426 48574
rect 263662 48338 299426 48574
rect 299662 48338 335426 48574
rect 335662 48338 371426 48574
rect 371662 48338 407426 48574
rect 407662 48338 443426 48574
rect 443662 48338 479426 48574
rect 479662 48338 515426 48574
rect 515662 48338 551426 48574
rect 551662 48338 591022 48574
rect 591258 48338 592350 48574
rect -8426 48326 592350 48338
rect -7506 48314 -6926 48326
rect 11254 48314 11834 48326
rect 47254 48314 47834 48326
rect 83254 48314 83834 48326
rect 119254 48314 119834 48326
rect 155254 48314 155834 48326
rect 191254 48314 191834 48326
rect 227254 48314 227834 48326
rect 263254 48314 263834 48326
rect 299254 48314 299834 48326
rect 335254 48314 335834 48326
rect 371254 48314 371834 48326
rect 407254 48314 407834 48326
rect 443254 48314 443834 48326
rect 479254 48314 479834 48326
rect 515254 48314 515834 48326
rect 551254 48314 551834 48326
rect 590850 48314 591430 48326
rect -5666 45426 -5086 45438
rect 7774 45426 8354 45438
rect 43774 45426 44354 45438
rect 79774 45426 80354 45438
rect 115774 45426 116354 45438
rect 151774 45426 152354 45438
rect 187774 45426 188354 45438
rect 223774 45426 224354 45438
rect 259774 45426 260354 45438
rect 295774 45426 296354 45438
rect 331774 45426 332354 45438
rect 367774 45426 368354 45438
rect 403774 45426 404354 45438
rect 439774 45426 440354 45438
rect 475774 45426 476354 45438
rect 511774 45426 512354 45438
rect 547774 45426 548354 45438
rect 589010 45426 589590 45438
rect -6586 45414 590510 45426
rect -6586 45178 -5494 45414
rect -5258 45178 7946 45414
rect 8182 45178 43946 45414
rect 44182 45178 79946 45414
rect 80182 45178 115946 45414
rect 116182 45178 151946 45414
rect 152182 45178 187946 45414
rect 188182 45178 223946 45414
rect 224182 45178 259946 45414
rect 260182 45178 295946 45414
rect 296182 45178 331946 45414
rect 332182 45178 367946 45414
rect 368182 45178 403946 45414
rect 404182 45178 439946 45414
rect 440182 45178 475946 45414
rect 476182 45178 511946 45414
rect 512182 45178 547946 45414
rect 548182 45178 589182 45414
rect 589418 45178 590510 45414
rect -6586 45094 590510 45178
rect -6586 44858 -5494 45094
rect -5258 44858 7946 45094
rect 8182 44858 43946 45094
rect 44182 44858 79946 45094
rect 80182 44858 115946 45094
rect 116182 44858 151946 45094
rect 152182 44858 187946 45094
rect 188182 44858 223946 45094
rect 224182 44858 259946 45094
rect 260182 44858 295946 45094
rect 296182 44858 331946 45094
rect 332182 44858 367946 45094
rect 368182 44858 403946 45094
rect 404182 44858 439946 45094
rect 440182 44858 475946 45094
rect 476182 44858 511946 45094
rect 512182 44858 547946 45094
rect 548182 44858 589182 45094
rect 589418 44858 590510 45094
rect -6586 44846 590510 44858
rect -5666 44834 -5086 44846
rect 7774 44834 8354 44846
rect 43774 44834 44354 44846
rect 79774 44834 80354 44846
rect 115774 44834 116354 44846
rect 151774 44834 152354 44846
rect 187774 44834 188354 44846
rect 223774 44834 224354 44846
rect 259774 44834 260354 44846
rect 295774 44834 296354 44846
rect 331774 44834 332354 44846
rect 367774 44834 368354 44846
rect 403774 44834 404354 44846
rect 439774 44834 440354 44846
rect 475774 44834 476354 44846
rect 511774 44834 512354 44846
rect 547774 44834 548354 44846
rect 589010 44834 589590 44846
rect -3826 41946 -3246 41958
rect 4294 41946 4874 41958
rect 40294 41946 40874 41958
rect 76294 41946 76874 41958
rect 112294 41946 112874 41958
rect 148294 41946 148874 41958
rect 184294 41946 184874 41958
rect 220294 41946 220874 41958
rect 256294 41946 256874 41958
rect 292294 41946 292874 41958
rect 328294 41946 328874 41958
rect 364294 41946 364874 41958
rect 400294 41946 400874 41958
rect 436294 41946 436874 41958
rect 472294 41946 472874 41958
rect 508294 41946 508874 41958
rect 544294 41946 544874 41958
rect 580294 41946 580874 41958
rect 587170 41946 587750 41958
rect -4746 41934 588670 41946
rect -4746 41698 -3654 41934
rect -3418 41698 4466 41934
rect 4702 41698 40466 41934
rect 40702 41698 76466 41934
rect 76702 41698 112466 41934
rect 112702 41698 148466 41934
rect 148702 41698 184466 41934
rect 184702 41698 220466 41934
rect 220702 41698 256466 41934
rect 256702 41698 292466 41934
rect 292702 41698 328466 41934
rect 328702 41698 364466 41934
rect 364702 41698 400466 41934
rect 400702 41698 436466 41934
rect 436702 41698 472466 41934
rect 472702 41698 508466 41934
rect 508702 41698 544466 41934
rect 544702 41698 580466 41934
rect 580702 41698 587342 41934
rect 587578 41698 588670 41934
rect -4746 41614 588670 41698
rect -4746 41378 -3654 41614
rect -3418 41378 4466 41614
rect 4702 41378 40466 41614
rect 40702 41378 76466 41614
rect 76702 41378 112466 41614
rect 112702 41378 148466 41614
rect 148702 41378 184466 41614
rect 184702 41378 220466 41614
rect 220702 41378 256466 41614
rect 256702 41378 292466 41614
rect 292702 41378 328466 41614
rect 328702 41378 364466 41614
rect 364702 41378 400466 41614
rect 400702 41378 436466 41614
rect 436702 41378 472466 41614
rect 472702 41378 508466 41614
rect 508702 41378 544466 41614
rect 544702 41378 580466 41614
rect 580702 41378 587342 41614
rect 587578 41378 588670 41614
rect -4746 41366 588670 41378
rect -3826 41354 -3246 41366
rect 4294 41354 4874 41366
rect 40294 41354 40874 41366
rect 76294 41354 76874 41366
rect 112294 41354 112874 41366
rect 148294 41354 148874 41366
rect 184294 41354 184874 41366
rect 220294 41354 220874 41366
rect 256294 41354 256874 41366
rect 292294 41354 292874 41366
rect 328294 41354 328874 41366
rect 364294 41354 364874 41366
rect 400294 41354 400874 41366
rect 436294 41354 436874 41366
rect 472294 41354 472874 41366
rect 508294 41354 508874 41366
rect 544294 41354 544874 41366
rect 580294 41354 580874 41366
rect 587170 41354 587750 41366
rect -1986 38466 -1406 38478
rect 814 38466 1394 38478
rect 36814 38466 37394 38478
rect 72814 38466 73394 38478
rect 108814 38466 109394 38478
rect 144814 38466 145394 38478
rect 180814 38466 181394 38478
rect 216814 38466 217394 38478
rect 252814 38466 253394 38478
rect 288814 38466 289394 38478
rect 324814 38466 325394 38478
rect 360814 38466 361394 38478
rect 396814 38466 397394 38478
rect 432814 38466 433394 38478
rect 468814 38466 469394 38478
rect 504814 38466 505394 38478
rect 540814 38466 541394 38478
rect 576814 38466 577394 38478
rect 585330 38466 585910 38478
rect -2906 38454 586830 38466
rect -2906 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586830 38454
rect -2906 38134 586830 38218
rect -2906 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586830 38134
rect -2906 37886 586830 37898
rect -1986 37874 -1406 37886
rect 814 37874 1394 37886
rect 36814 37874 37394 37886
rect 72814 37874 73394 37886
rect 108814 37874 109394 37886
rect 144814 37874 145394 37886
rect 180814 37874 181394 37886
rect 216814 37874 217394 37886
rect 252814 37874 253394 37886
rect 288814 37874 289394 37886
rect 324814 37874 325394 37886
rect 360814 37874 361394 37886
rect 396814 37874 397394 37886
rect 432814 37874 433394 37886
rect 468814 37874 469394 37886
rect 504814 37874 505394 37886
rect 540814 37874 541394 37886
rect 576814 37874 577394 37886
rect 585330 37874 585910 37886
rect -8426 30906 -7846 30918
rect 29254 30906 29834 30918
rect 65254 30906 65834 30918
rect 101254 30906 101834 30918
rect 137254 30906 137834 30918
rect 173254 30906 173834 30918
rect 209254 30906 209834 30918
rect 245254 30906 245834 30918
rect 281254 30906 281834 30918
rect 317254 30906 317834 30918
rect 353254 30906 353834 30918
rect 389254 30906 389834 30918
rect 425254 30906 425834 30918
rect 461254 30906 461834 30918
rect 497254 30906 497834 30918
rect 533254 30906 533834 30918
rect 569254 30906 569834 30918
rect 591770 30906 592350 30918
rect -8426 30894 592350 30906
rect -8426 30658 -8254 30894
rect -8018 30658 29426 30894
rect 29662 30658 65426 30894
rect 65662 30658 101426 30894
rect 101662 30658 137426 30894
rect 137662 30658 173426 30894
rect 173662 30658 209426 30894
rect 209662 30658 245426 30894
rect 245662 30658 281426 30894
rect 281662 30658 317426 30894
rect 317662 30658 353426 30894
rect 353662 30658 389426 30894
rect 389662 30658 425426 30894
rect 425662 30658 461426 30894
rect 461662 30658 497426 30894
rect 497662 30658 533426 30894
rect 533662 30658 569426 30894
rect 569662 30658 591942 30894
rect 592178 30658 592350 30894
rect -8426 30574 592350 30658
rect -8426 30338 -8254 30574
rect -8018 30338 29426 30574
rect 29662 30338 65426 30574
rect 65662 30338 101426 30574
rect 101662 30338 137426 30574
rect 137662 30338 173426 30574
rect 173662 30338 209426 30574
rect 209662 30338 245426 30574
rect 245662 30338 281426 30574
rect 281662 30338 317426 30574
rect 317662 30338 353426 30574
rect 353662 30338 389426 30574
rect 389662 30338 425426 30574
rect 425662 30338 461426 30574
rect 461662 30338 497426 30574
rect 497662 30338 533426 30574
rect 533662 30338 569426 30574
rect 569662 30338 591942 30574
rect 592178 30338 592350 30574
rect -8426 30326 592350 30338
rect -8426 30314 -7846 30326
rect 29254 30314 29834 30326
rect 65254 30314 65834 30326
rect 101254 30314 101834 30326
rect 137254 30314 137834 30326
rect 173254 30314 173834 30326
rect 209254 30314 209834 30326
rect 245254 30314 245834 30326
rect 281254 30314 281834 30326
rect 317254 30314 317834 30326
rect 353254 30314 353834 30326
rect 389254 30314 389834 30326
rect 425254 30314 425834 30326
rect 461254 30314 461834 30326
rect 497254 30314 497834 30326
rect 533254 30314 533834 30326
rect 569254 30314 569834 30326
rect 591770 30314 592350 30326
rect -6586 27426 -6006 27438
rect 25774 27426 26354 27438
rect 61774 27426 62354 27438
rect 97774 27426 98354 27438
rect 133774 27426 134354 27438
rect 169774 27426 170354 27438
rect 205774 27426 206354 27438
rect 241774 27426 242354 27438
rect 277774 27426 278354 27438
rect 313774 27426 314354 27438
rect 349774 27426 350354 27438
rect 385774 27426 386354 27438
rect 421774 27426 422354 27438
rect 457774 27426 458354 27438
rect 493774 27426 494354 27438
rect 529774 27426 530354 27438
rect 565774 27426 566354 27438
rect 589930 27426 590510 27438
rect -6586 27414 590510 27426
rect -6586 27178 -6414 27414
rect -6178 27178 25946 27414
rect 26182 27178 61946 27414
rect 62182 27178 97946 27414
rect 98182 27178 133946 27414
rect 134182 27178 169946 27414
rect 170182 27178 205946 27414
rect 206182 27178 241946 27414
rect 242182 27178 277946 27414
rect 278182 27178 313946 27414
rect 314182 27178 349946 27414
rect 350182 27178 385946 27414
rect 386182 27178 421946 27414
rect 422182 27178 457946 27414
rect 458182 27178 493946 27414
rect 494182 27178 529946 27414
rect 530182 27178 565946 27414
rect 566182 27178 590102 27414
rect 590338 27178 590510 27414
rect -6586 27094 590510 27178
rect -6586 26858 -6414 27094
rect -6178 26858 25946 27094
rect 26182 26858 61946 27094
rect 62182 26858 97946 27094
rect 98182 26858 133946 27094
rect 134182 26858 169946 27094
rect 170182 26858 205946 27094
rect 206182 26858 241946 27094
rect 242182 26858 277946 27094
rect 278182 26858 313946 27094
rect 314182 26858 349946 27094
rect 350182 26858 385946 27094
rect 386182 26858 421946 27094
rect 422182 26858 457946 27094
rect 458182 26858 493946 27094
rect 494182 26858 529946 27094
rect 530182 26858 565946 27094
rect 566182 26858 590102 27094
rect 590338 26858 590510 27094
rect -6586 26846 590510 26858
rect -6586 26834 -6006 26846
rect 25774 26834 26354 26846
rect 61774 26834 62354 26846
rect 97774 26834 98354 26846
rect 133774 26834 134354 26846
rect 169774 26834 170354 26846
rect 205774 26834 206354 26846
rect 241774 26834 242354 26846
rect 277774 26834 278354 26846
rect 313774 26834 314354 26846
rect 349774 26834 350354 26846
rect 385774 26834 386354 26846
rect 421774 26834 422354 26846
rect 457774 26834 458354 26846
rect 493774 26834 494354 26846
rect 529774 26834 530354 26846
rect 565774 26834 566354 26846
rect 589930 26834 590510 26846
rect -4746 23946 -4166 23958
rect 22294 23946 22874 23958
rect 58294 23946 58874 23958
rect 94294 23946 94874 23958
rect 130294 23946 130874 23958
rect 166294 23946 166874 23958
rect 202294 23946 202874 23958
rect 238294 23946 238874 23958
rect 274294 23946 274874 23958
rect 310294 23946 310874 23958
rect 346294 23946 346874 23958
rect 382294 23946 382874 23958
rect 418294 23946 418874 23958
rect 454294 23946 454874 23958
rect 490294 23946 490874 23958
rect 526294 23946 526874 23958
rect 562294 23946 562874 23958
rect 588090 23946 588670 23958
rect -4746 23934 588670 23946
rect -4746 23698 -4574 23934
rect -4338 23698 22466 23934
rect 22702 23698 58466 23934
rect 58702 23698 94466 23934
rect 94702 23698 130466 23934
rect 130702 23698 166466 23934
rect 166702 23698 202466 23934
rect 202702 23698 238466 23934
rect 238702 23698 274466 23934
rect 274702 23698 310466 23934
rect 310702 23698 346466 23934
rect 346702 23698 382466 23934
rect 382702 23698 418466 23934
rect 418702 23698 454466 23934
rect 454702 23698 490466 23934
rect 490702 23698 526466 23934
rect 526702 23698 562466 23934
rect 562702 23698 588262 23934
rect 588498 23698 588670 23934
rect -4746 23614 588670 23698
rect -4746 23378 -4574 23614
rect -4338 23378 22466 23614
rect 22702 23378 58466 23614
rect 58702 23378 94466 23614
rect 94702 23378 130466 23614
rect 130702 23378 166466 23614
rect 166702 23378 202466 23614
rect 202702 23378 238466 23614
rect 238702 23378 274466 23614
rect 274702 23378 310466 23614
rect 310702 23378 346466 23614
rect 346702 23378 382466 23614
rect 382702 23378 418466 23614
rect 418702 23378 454466 23614
rect 454702 23378 490466 23614
rect 490702 23378 526466 23614
rect 526702 23378 562466 23614
rect 562702 23378 588262 23614
rect 588498 23378 588670 23614
rect -4746 23366 588670 23378
rect -4746 23354 -4166 23366
rect 22294 23354 22874 23366
rect 58294 23354 58874 23366
rect 94294 23354 94874 23366
rect 130294 23354 130874 23366
rect 166294 23354 166874 23366
rect 202294 23354 202874 23366
rect 238294 23354 238874 23366
rect 274294 23354 274874 23366
rect 310294 23354 310874 23366
rect 346294 23354 346874 23366
rect 382294 23354 382874 23366
rect 418294 23354 418874 23366
rect 454294 23354 454874 23366
rect 490294 23354 490874 23366
rect 526294 23354 526874 23366
rect 562294 23354 562874 23366
rect 588090 23354 588670 23366
rect -2906 20466 -2326 20478
rect 18814 20466 19394 20478
rect 54814 20466 55394 20478
rect 90814 20466 91394 20478
rect 126814 20466 127394 20478
rect 162814 20466 163394 20478
rect 198814 20466 199394 20478
rect 234814 20466 235394 20478
rect 270814 20466 271394 20478
rect 306814 20466 307394 20478
rect 342814 20466 343394 20478
rect 378814 20466 379394 20478
rect 414814 20466 415394 20478
rect 450814 20466 451394 20478
rect 486814 20466 487394 20478
rect 522814 20466 523394 20478
rect 558814 20466 559394 20478
rect 586250 20466 586830 20478
rect -2906 20454 586830 20466
rect -2906 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586830 20454
rect -2906 20134 586830 20218
rect -2906 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586830 20134
rect -2906 19886 586830 19898
rect -2906 19874 -2326 19886
rect 18814 19874 19394 19886
rect 54814 19874 55394 19886
rect 90814 19874 91394 19886
rect 126814 19874 127394 19886
rect 162814 19874 163394 19886
rect 198814 19874 199394 19886
rect 234814 19874 235394 19886
rect 270814 19874 271394 19886
rect 306814 19874 307394 19886
rect 342814 19874 343394 19886
rect 378814 19874 379394 19886
rect 414814 19874 415394 19886
rect 450814 19874 451394 19886
rect 486814 19874 487394 19886
rect 522814 19874 523394 19886
rect 558814 19874 559394 19886
rect 586250 19874 586830 19886
rect -7506 12906 -6926 12918
rect 11254 12906 11834 12918
rect 47254 12906 47834 12918
rect 83254 12906 83834 12918
rect 119254 12906 119834 12918
rect 155254 12906 155834 12918
rect 191254 12906 191834 12918
rect 227254 12906 227834 12918
rect 263254 12906 263834 12918
rect 299254 12906 299834 12918
rect 335254 12906 335834 12918
rect 371254 12906 371834 12918
rect 407254 12906 407834 12918
rect 443254 12906 443834 12918
rect 479254 12906 479834 12918
rect 515254 12906 515834 12918
rect 551254 12906 551834 12918
rect 590850 12906 591430 12918
rect -8426 12894 592350 12906
rect -8426 12658 -7334 12894
rect -7098 12658 11426 12894
rect 11662 12658 47426 12894
rect 47662 12658 83426 12894
rect 83662 12658 119426 12894
rect 119662 12658 155426 12894
rect 155662 12658 191426 12894
rect 191662 12658 227426 12894
rect 227662 12658 263426 12894
rect 263662 12658 299426 12894
rect 299662 12658 335426 12894
rect 335662 12658 371426 12894
rect 371662 12658 407426 12894
rect 407662 12658 443426 12894
rect 443662 12658 479426 12894
rect 479662 12658 515426 12894
rect 515662 12658 551426 12894
rect 551662 12658 591022 12894
rect 591258 12658 592350 12894
rect -8426 12574 592350 12658
rect -8426 12338 -7334 12574
rect -7098 12338 11426 12574
rect 11662 12338 47426 12574
rect 47662 12338 83426 12574
rect 83662 12338 119426 12574
rect 119662 12338 155426 12574
rect 155662 12338 191426 12574
rect 191662 12338 227426 12574
rect 227662 12338 263426 12574
rect 263662 12338 299426 12574
rect 299662 12338 335426 12574
rect 335662 12338 371426 12574
rect 371662 12338 407426 12574
rect 407662 12338 443426 12574
rect 443662 12338 479426 12574
rect 479662 12338 515426 12574
rect 515662 12338 551426 12574
rect 551662 12338 591022 12574
rect 591258 12338 592350 12574
rect -8426 12326 592350 12338
rect -7506 12314 -6926 12326
rect 11254 12314 11834 12326
rect 47254 12314 47834 12326
rect 83254 12314 83834 12326
rect 119254 12314 119834 12326
rect 155254 12314 155834 12326
rect 191254 12314 191834 12326
rect 227254 12314 227834 12326
rect 263254 12314 263834 12326
rect 299254 12314 299834 12326
rect 335254 12314 335834 12326
rect 371254 12314 371834 12326
rect 407254 12314 407834 12326
rect 443254 12314 443834 12326
rect 479254 12314 479834 12326
rect 515254 12314 515834 12326
rect 551254 12314 551834 12326
rect 590850 12314 591430 12326
rect -5666 9426 -5086 9438
rect 7774 9426 8354 9438
rect 43774 9426 44354 9438
rect 79774 9426 80354 9438
rect 115774 9426 116354 9438
rect 151774 9426 152354 9438
rect 187774 9426 188354 9438
rect 223774 9426 224354 9438
rect 259774 9426 260354 9438
rect 295774 9426 296354 9438
rect 331774 9426 332354 9438
rect 367774 9426 368354 9438
rect 403774 9426 404354 9438
rect 439774 9426 440354 9438
rect 475774 9426 476354 9438
rect 511774 9426 512354 9438
rect 547774 9426 548354 9438
rect 589010 9426 589590 9438
rect -6586 9414 590510 9426
rect -6586 9178 -5494 9414
rect -5258 9178 7946 9414
rect 8182 9178 43946 9414
rect 44182 9178 79946 9414
rect 80182 9178 115946 9414
rect 116182 9178 151946 9414
rect 152182 9178 187946 9414
rect 188182 9178 223946 9414
rect 224182 9178 259946 9414
rect 260182 9178 295946 9414
rect 296182 9178 331946 9414
rect 332182 9178 367946 9414
rect 368182 9178 403946 9414
rect 404182 9178 439946 9414
rect 440182 9178 475946 9414
rect 476182 9178 511946 9414
rect 512182 9178 547946 9414
rect 548182 9178 589182 9414
rect 589418 9178 590510 9414
rect -6586 9094 590510 9178
rect -6586 8858 -5494 9094
rect -5258 8858 7946 9094
rect 8182 8858 43946 9094
rect 44182 8858 79946 9094
rect 80182 8858 115946 9094
rect 116182 8858 151946 9094
rect 152182 8858 187946 9094
rect 188182 8858 223946 9094
rect 224182 8858 259946 9094
rect 260182 8858 295946 9094
rect 296182 8858 331946 9094
rect 332182 8858 367946 9094
rect 368182 8858 403946 9094
rect 404182 8858 439946 9094
rect 440182 8858 475946 9094
rect 476182 8858 511946 9094
rect 512182 8858 547946 9094
rect 548182 8858 589182 9094
rect 589418 8858 590510 9094
rect -6586 8846 590510 8858
rect -5666 8834 -5086 8846
rect 7774 8834 8354 8846
rect 43774 8834 44354 8846
rect 79774 8834 80354 8846
rect 115774 8834 116354 8846
rect 151774 8834 152354 8846
rect 187774 8834 188354 8846
rect 223774 8834 224354 8846
rect 259774 8834 260354 8846
rect 295774 8834 296354 8846
rect 331774 8834 332354 8846
rect 367774 8834 368354 8846
rect 403774 8834 404354 8846
rect 439774 8834 440354 8846
rect 475774 8834 476354 8846
rect 511774 8834 512354 8846
rect 547774 8834 548354 8846
rect 589010 8834 589590 8846
rect -3826 5946 -3246 5958
rect 4294 5946 4874 5958
rect 40294 5946 40874 5958
rect 76294 5946 76874 5958
rect 112294 5946 112874 5958
rect 148294 5946 148874 5958
rect 184294 5946 184874 5958
rect 220294 5946 220874 5958
rect 256294 5946 256874 5958
rect 292294 5946 292874 5958
rect 328294 5946 328874 5958
rect 364294 5946 364874 5958
rect 400294 5946 400874 5958
rect 436294 5946 436874 5958
rect 472294 5946 472874 5958
rect 508294 5946 508874 5958
rect 544294 5946 544874 5958
rect 580294 5946 580874 5958
rect 587170 5946 587750 5958
rect -4746 5934 588670 5946
rect -4746 5698 -3654 5934
rect -3418 5698 4466 5934
rect 4702 5698 40466 5934
rect 40702 5698 76466 5934
rect 76702 5698 112466 5934
rect 112702 5698 148466 5934
rect 148702 5698 184466 5934
rect 184702 5698 220466 5934
rect 220702 5698 256466 5934
rect 256702 5698 292466 5934
rect 292702 5698 328466 5934
rect 328702 5698 364466 5934
rect 364702 5698 400466 5934
rect 400702 5698 436466 5934
rect 436702 5698 472466 5934
rect 472702 5698 508466 5934
rect 508702 5698 544466 5934
rect 544702 5698 580466 5934
rect 580702 5698 587342 5934
rect 587578 5698 588670 5934
rect -4746 5614 588670 5698
rect -4746 5378 -3654 5614
rect -3418 5378 4466 5614
rect 4702 5378 40466 5614
rect 40702 5378 76466 5614
rect 76702 5378 112466 5614
rect 112702 5378 148466 5614
rect 148702 5378 184466 5614
rect 184702 5378 220466 5614
rect 220702 5378 256466 5614
rect 256702 5378 292466 5614
rect 292702 5378 328466 5614
rect 328702 5378 364466 5614
rect 364702 5378 400466 5614
rect 400702 5378 436466 5614
rect 436702 5378 472466 5614
rect 472702 5378 508466 5614
rect 508702 5378 544466 5614
rect 544702 5378 580466 5614
rect 580702 5378 587342 5614
rect 587578 5378 588670 5614
rect -4746 5366 588670 5378
rect -3826 5354 -3246 5366
rect 4294 5354 4874 5366
rect 40294 5354 40874 5366
rect 76294 5354 76874 5366
rect 112294 5354 112874 5366
rect 148294 5354 148874 5366
rect 184294 5354 184874 5366
rect 220294 5354 220874 5366
rect 256294 5354 256874 5366
rect 292294 5354 292874 5366
rect 328294 5354 328874 5366
rect 364294 5354 364874 5366
rect 400294 5354 400874 5366
rect 436294 5354 436874 5366
rect 472294 5354 472874 5366
rect 508294 5354 508874 5366
rect 544294 5354 544874 5366
rect 580294 5354 580874 5366
rect 587170 5354 587750 5366
rect -1986 2466 -1406 2478
rect 814 2466 1394 2478
rect 36814 2466 37394 2478
rect 72814 2466 73394 2478
rect 108814 2466 109394 2478
rect 144814 2466 145394 2478
rect 180814 2466 181394 2478
rect 216814 2466 217394 2478
rect 252814 2466 253394 2478
rect 288814 2466 289394 2478
rect 324814 2466 325394 2478
rect 360814 2466 361394 2478
rect 396814 2466 397394 2478
rect 432814 2466 433394 2478
rect 468814 2466 469394 2478
rect 504814 2466 505394 2478
rect 540814 2466 541394 2478
rect 576814 2466 577394 2478
rect 585330 2466 585910 2478
rect -2906 2454 586830 2466
rect -2906 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586830 2454
rect -2906 2134 586830 2218
rect -2906 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586830 2134
rect -2906 1886 586830 1898
rect -1986 1874 -1406 1886
rect 814 1874 1394 1886
rect 36814 1874 37394 1886
rect 72814 1874 73394 1886
rect 108814 1874 109394 1886
rect 144814 1874 145394 1886
rect 180814 1874 181394 1886
rect 216814 1874 217394 1886
rect 252814 1874 253394 1886
rect 288814 1874 289394 1886
rect 324814 1874 325394 1886
rect 360814 1874 361394 1886
rect 396814 1874 397394 1886
rect 432814 1874 433394 1886
rect 468814 1874 469394 1886
rect 504814 1874 505394 1886
rect 540814 1874 541394 1886
rect 576814 1874 577394 1886
rect 585330 1874 585910 1886
rect -1986 -334 -1406 -322
rect 814 -334 1394 -322
rect 36814 -334 37394 -322
rect 72814 -334 73394 -322
rect 108814 -334 109394 -322
rect 144814 -334 145394 -322
rect 180814 -334 181394 -322
rect 216814 -334 217394 -322
rect 252814 -334 253394 -322
rect 288814 -334 289394 -322
rect 324814 -334 325394 -322
rect 360814 -334 361394 -322
rect 396814 -334 397394 -322
rect 432814 -334 433394 -322
rect 468814 -334 469394 -322
rect 504814 -334 505394 -322
rect 540814 -334 541394 -322
rect 576814 -334 577394 -322
rect 585330 -334 585910 -322
rect -1986 -346 585910 -334
rect -1986 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585910 -346
rect -1986 -666 585910 -582
rect -1986 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585910 -666
rect -1986 -914 585910 -902
rect -1986 -926 -1406 -914
rect 814 -926 1394 -914
rect 36814 -926 37394 -914
rect 72814 -926 73394 -914
rect 108814 -926 109394 -914
rect 144814 -926 145394 -914
rect 180814 -926 181394 -914
rect 216814 -926 217394 -914
rect 252814 -926 253394 -914
rect 288814 -926 289394 -914
rect 324814 -926 325394 -914
rect 360814 -926 361394 -914
rect 396814 -926 397394 -914
rect 432814 -926 433394 -914
rect 468814 -926 469394 -914
rect 504814 -926 505394 -914
rect 540814 -926 541394 -914
rect 576814 -926 577394 -914
rect 585330 -926 585910 -914
rect -2906 -1254 -2326 -1242
rect 18814 -1254 19394 -1242
rect 54814 -1254 55394 -1242
rect 90814 -1254 91394 -1242
rect 126814 -1254 127394 -1242
rect 162814 -1254 163394 -1242
rect 198814 -1254 199394 -1242
rect 234814 -1254 235394 -1242
rect 270814 -1254 271394 -1242
rect 306814 -1254 307394 -1242
rect 342814 -1254 343394 -1242
rect 378814 -1254 379394 -1242
rect 414814 -1254 415394 -1242
rect 450814 -1254 451394 -1242
rect 486814 -1254 487394 -1242
rect 522814 -1254 523394 -1242
rect 558814 -1254 559394 -1242
rect 586250 -1254 586830 -1242
rect -2906 -1266 586830 -1254
rect -2906 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586830 -1266
rect -2906 -1586 586830 -1502
rect -2906 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586830 -1586
rect -2906 -1834 586830 -1822
rect -2906 -1846 -2326 -1834
rect 18814 -1846 19394 -1834
rect 54814 -1846 55394 -1834
rect 90814 -1846 91394 -1834
rect 126814 -1846 127394 -1834
rect 162814 -1846 163394 -1834
rect 198814 -1846 199394 -1834
rect 234814 -1846 235394 -1834
rect 270814 -1846 271394 -1834
rect 306814 -1846 307394 -1834
rect 342814 -1846 343394 -1834
rect 378814 -1846 379394 -1834
rect 414814 -1846 415394 -1834
rect 450814 -1846 451394 -1834
rect 486814 -1846 487394 -1834
rect 522814 -1846 523394 -1834
rect 558814 -1846 559394 -1834
rect 586250 -1846 586830 -1834
rect -3826 -2174 -3246 -2162
rect 4294 -2174 4874 -2162
rect 40294 -2174 40874 -2162
rect 76294 -2174 76874 -2162
rect 112294 -2174 112874 -2162
rect 148294 -2174 148874 -2162
rect 184294 -2174 184874 -2162
rect 220294 -2174 220874 -2162
rect 256294 -2174 256874 -2162
rect 292294 -2174 292874 -2162
rect 328294 -2174 328874 -2162
rect 364294 -2174 364874 -2162
rect 400294 -2174 400874 -2162
rect 436294 -2174 436874 -2162
rect 472294 -2174 472874 -2162
rect 508294 -2174 508874 -2162
rect 544294 -2174 544874 -2162
rect 580294 -2174 580874 -2162
rect 587170 -2174 587750 -2162
rect -3826 -2186 587750 -2174
rect -3826 -2422 -3654 -2186
rect -3418 -2422 4466 -2186
rect 4702 -2422 40466 -2186
rect 40702 -2422 76466 -2186
rect 76702 -2422 112466 -2186
rect 112702 -2422 148466 -2186
rect 148702 -2422 184466 -2186
rect 184702 -2422 220466 -2186
rect 220702 -2422 256466 -2186
rect 256702 -2422 292466 -2186
rect 292702 -2422 328466 -2186
rect 328702 -2422 364466 -2186
rect 364702 -2422 400466 -2186
rect 400702 -2422 436466 -2186
rect 436702 -2422 472466 -2186
rect 472702 -2422 508466 -2186
rect 508702 -2422 544466 -2186
rect 544702 -2422 580466 -2186
rect 580702 -2422 587342 -2186
rect 587578 -2422 587750 -2186
rect -3826 -2506 587750 -2422
rect -3826 -2742 -3654 -2506
rect -3418 -2742 4466 -2506
rect 4702 -2742 40466 -2506
rect 40702 -2742 76466 -2506
rect 76702 -2742 112466 -2506
rect 112702 -2742 148466 -2506
rect 148702 -2742 184466 -2506
rect 184702 -2742 220466 -2506
rect 220702 -2742 256466 -2506
rect 256702 -2742 292466 -2506
rect 292702 -2742 328466 -2506
rect 328702 -2742 364466 -2506
rect 364702 -2742 400466 -2506
rect 400702 -2742 436466 -2506
rect 436702 -2742 472466 -2506
rect 472702 -2742 508466 -2506
rect 508702 -2742 544466 -2506
rect 544702 -2742 580466 -2506
rect 580702 -2742 587342 -2506
rect 587578 -2742 587750 -2506
rect -3826 -2754 587750 -2742
rect -3826 -2766 -3246 -2754
rect 4294 -2766 4874 -2754
rect 40294 -2766 40874 -2754
rect 76294 -2766 76874 -2754
rect 112294 -2766 112874 -2754
rect 148294 -2766 148874 -2754
rect 184294 -2766 184874 -2754
rect 220294 -2766 220874 -2754
rect 256294 -2766 256874 -2754
rect 292294 -2766 292874 -2754
rect 328294 -2766 328874 -2754
rect 364294 -2766 364874 -2754
rect 400294 -2766 400874 -2754
rect 436294 -2766 436874 -2754
rect 472294 -2766 472874 -2754
rect 508294 -2766 508874 -2754
rect 544294 -2766 544874 -2754
rect 580294 -2766 580874 -2754
rect 587170 -2766 587750 -2754
rect -4746 -3094 -4166 -3082
rect 22294 -3094 22874 -3082
rect 58294 -3094 58874 -3082
rect 94294 -3094 94874 -3082
rect 130294 -3094 130874 -3082
rect 166294 -3094 166874 -3082
rect 202294 -3094 202874 -3082
rect 238294 -3094 238874 -3082
rect 274294 -3094 274874 -3082
rect 310294 -3094 310874 -3082
rect 346294 -3094 346874 -3082
rect 382294 -3094 382874 -3082
rect 418294 -3094 418874 -3082
rect 454294 -3094 454874 -3082
rect 490294 -3094 490874 -3082
rect 526294 -3094 526874 -3082
rect 562294 -3094 562874 -3082
rect 588090 -3094 588670 -3082
rect -4746 -3106 588670 -3094
rect -4746 -3342 -4574 -3106
rect -4338 -3342 22466 -3106
rect 22702 -3342 58466 -3106
rect 58702 -3342 94466 -3106
rect 94702 -3342 130466 -3106
rect 130702 -3342 166466 -3106
rect 166702 -3342 202466 -3106
rect 202702 -3342 238466 -3106
rect 238702 -3342 274466 -3106
rect 274702 -3342 310466 -3106
rect 310702 -3342 346466 -3106
rect 346702 -3342 382466 -3106
rect 382702 -3342 418466 -3106
rect 418702 -3342 454466 -3106
rect 454702 -3342 490466 -3106
rect 490702 -3342 526466 -3106
rect 526702 -3342 562466 -3106
rect 562702 -3342 588262 -3106
rect 588498 -3342 588670 -3106
rect -4746 -3426 588670 -3342
rect -4746 -3662 -4574 -3426
rect -4338 -3662 22466 -3426
rect 22702 -3662 58466 -3426
rect 58702 -3662 94466 -3426
rect 94702 -3662 130466 -3426
rect 130702 -3662 166466 -3426
rect 166702 -3662 202466 -3426
rect 202702 -3662 238466 -3426
rect 238702 -3662 274466 -3426
rect 274702 -3662 310466 -3426
rect 310702 -3662 346466 -3426
rect 346702 -3662 382466 -3426
rect 382702 -3662 418466 -3426
rect 418702 -3662 454466 -3426
rect 454702 -3662 490466 -3426
rect 490702 -3662 526466 -3426
rect 526702 -3662 562466 -3426
rect 562702 -3662 588262 -3426
rect 588498 -3662 588670 -3426
rect -4746 -3674 588670 -3662
rect -4746 -3686 -4166 -3674
rect 22294 -3686 22874 -3674
rect 58294 -3686 58874 -3674
rect 94294 -3686 94874 -3674
rect 130294 -3686 130874 -3674
rect 166294 -3686 166874 -3674
rect 202294 -3686 202874 -3674
rect 238294 -3686 238874 -3674
rect 274294 -3686 274874 -3674
rect 310294 -3686 310874 -3674
rect 346294 -3686 346874 -3674
rect 382294 -3686 382874 -3674
rect 418294 -3686 418874 -3674
rect 454294 -3686 454874 -3674
rect 490294 -3686 490874 -3674
rect 526294 -3686 526874 -3674
rect 562294 -3686 562874 -3674
rect 588090 -3686 588670 -3674
rect -5666 -4014 -5086 -4002
rect 7774 -4014 8354 -4002
rect 43774 -4014 44354 -4002
rect 79774 -4014 80354 -4002
rect 115774 -4014 116354 -4002
rect 151774 -4014 152354 -4002
rect 187774 -4014 188354 -4002
rect 223774 -4014 224354 -4002
rect 259774 -4014 260354 -4002
rect 295774 -4014 296354 -4002
rect 331774 -4014 332354 -4002
rect 367774 -4014 368354 -4002
rect 403774 -4014 404354 -4002
rect 439774 -4014 440354 -4002
rect 475774 -4014 476354 -4002
rect 511774 -4014 512354 -4002
rect 547774 -4014 548354 -4002
rect 589010 -4014 589590 -4002
rect -5666 -4026 589590 -4014
rect -5666 -4262 -5494 -4026
rect -5258 -4262 7946 -4026
rect 8182 -4262 43946 -4026
rect 44182 -4262 79946 -4026
rect 80182 -4262 115946 -4026
rect 116182 -4262 151946 -4026
rect 152182 -4262 187946 -4026
rect 188182 -4262 223946 -4026
rect 224182 -4262 259946 -4026
rect 260182 -4262 295946 -4026
rect 296182 -4262 331946 -4026
rect 332182 -4262 367946 -4026
rect 368182 -4262 403946 -4026
rect 404182 -4262 439946 -4026
rect 440182 -4262 475946 -4026
rect 476182 -4262 511946 -4026
rect 512182 -4262 547946 -4026
rect 548182 -4262 589182 -4026
rect 589418 -4262 589590 -4026
rect -5666 -4346 589590 -4262
rect -5666 -4582 -5494 -4346
rect -5258 -4582 7946 -4346
rect 8182 -4582 43946 -4346
rect 44182 -4582 79946 -4346
rect 80182 -4582 115946 -4346
rect 116182 -4582 151946 -4346
rect 152182 -4582 187946 -4346
rect 188182 -4582 223946 -4346
rect 224182 -4582 259946 -4346
rect 260182 -4582 295946 -4346
rect 296182 -4582 331946 -4346
rect 332182 -4582 367946 -4346
rect 368182 -4582 403946 -4346
rect 404182 -4582 439946 -4346
rect 440182 -4582 475946 -4346
rect 476182 -4582 511946 -4346
rect 512182 -4582 547946 -4346
rect 548182 -4582 589182 -4346
rect 589418 -4582 589590 -4346
rect -5666 -4594 589590 -4582
rect -5666 -4606 -5086 -4594
rect 7774 -4606 8354 -4594
rect 43774 -4606 44354 -4594
rect 79774 -4606 80354 -4594
rect 115774 -4606 116354 -4594
rect 151774 -4606 152354 -4594
rect 187774 -4606 188354 -4594
rect 223774 -4606 224354 -4594
rect 259774 -4606 260354 -4594
rect 295774 -4606 296354 -4594
rect 331774 -4606 332354 -4594
rect 367774 -4606 368354 -4594
rect 403774 -4606 404354 -4594
rect 439774 -4606 440354 -4594
rect 475774 -4606 476354 -4594
rect 511774 -4606 512354 -4594
rect 547774 -4606 548354 -4594
rect 589010 -4606 589590 -4594
rect -6586 -4934 -6006 -4922
rect 25774 -4934 26354 -4922
rect 61774 -4934 62354 -4922
rect 97774 -4934 98354 -4922
rect 133774 -4934 134354 -4922
rect 169774 -4934 170354 -4922
rect 205774 -4934 206354 -4922
rect 241774 -4934 242354 -4922
rect 277774 -4934 278354 -4922
rect 313774 -4934 314354 -4922
rect 349774 -4934 350354 -4922
rect 385774 -4934 386354 -4922
rect 421774 -4934 422354 -4922
rect 457774 -4934 458354 -4922
rect 493774 -4934 494354 -4922
rect 529774 -4934 530354 -4922
rect 565774 -4934 566354 -4922
rect 589930 -4934 590510 -4922
rect -6586 -4946 590510 -4934
rect -6586 -5182 -6414 -4946
rect -6178 -5182 25946 -4946
rect 26182 -5182 61946 -4946
rect 62182 -5182 97946 -4946
rect 98182 -5182 133946 -4946
rect 134182 -5182 169946 -4946
rect 170182 -5182 205946 -4946
rect 206182 -5182 241946 -4946
rect 242182 -5182 277946 -4946
rect 278182 -5182 313946 -4946
rect 314182 -5182 349946 -4946
rect 350182 -5182 385946 -4946
rect 386182 -5182 421946 -4946
rect 422182 -5182 457946 -4946
rect 458182 -5182 493946 -4946
rect 494182 -5182 529946 -4946
rect 530182 -5182 565946 -4946
rect 566182 -5182 590102 -4946
rect 590338 -5182 590510 -4946
rect -6586 -5266 590510 -5182
rect -6586 -5502 -6414 -5266
rect -6178 -5502 25946 -5266
rect 26182 -5502 61946 -5266
rect 62182 -5502 97946 -5266
rect 98182 -5502 133946 -5266
rect 134182 -5502 169946 -5266
rect 170182 -5502 205946 -5266
rect 206182 -5502 241946 -5266
rect 242182 -5502 277946 -5266
rect 278182 -5502 313946 -5266
rect 314182 -5502 349946 -5266
rect 350182 -5502 385946 -5266
rect 386182 -5502 421946 -5266
rect 422182 -5502 457946 -5266
rect 458182 -5502 493946 -5266
rect 494182 -5502 529946 -5266
rect 530182 -5502 565946 -5266
rect 566182 -5502 590102 -5266
rect 590338 -5502 590510 -5266
rect -6586 -5514 590510 -5502
rect -6586 -5526 -6006 -5514
rect 25774 -5526 26354 -5514
rect 61774 -5526 62354 -5514
rect 97774 -5526 98354 -5514
rect 133774 -5526 134354 -5514
rect 169774 -5526 170354 -5514
rect 205774 -5526 206354 -5514
rect 241774 -5526 242354 -5514
rect 277774 -5526 278354 -5514
rect 313774 -5526 314354 -5514
rect 349774 -5526 350354 -5514
rect 385774 -5526 386354 -5514
rect 421774 -5526 422354 -5514
rect 457774 -5526 458354 -5514
rect 493774 -5526 494354 -5514
rect 529774 -5526 530354 -5514
rect 565774 -5526 566354 -5514
rect 589930 -5526 590510 -5514
rect -7506 -5854 -6926 -5842
rect 11254 -5854 11834 -5842
rect 47254 -5854 47834 -5842
rect 83254 -5854 83834 -5842
rect 119254 -5854 119834 -5842
rect 155254 -5854 155834 -5842
rect 191254 -5854 191834 -5842
rect 227254 -5854 227834 -5842
rect 263254 -5854 263834 -5842
rect 299254 -5854 299834 -5842
rect 335254 -5854 335834 -5842
rect 371254 -5854 371834 -5842
rect 407254 -5854 407834 -5842
rect 443254 -5854 443834 -5842
rect 479254 -5854 479834 -5842
rect 515254 -5854 515834 -5842
rect 551254 -5854 551834 -5842
rect 590850 -5854 591430 -5842
rect -7506 -5866 591430 -5854
rect -7506 -6102 -7334 -5866
rect -7098 -6102 11426 -5866
rect 11662 -6102 47426 -5866
rect 47662 -6102 83426 -5866
rect 83662 -6102 119426 -5866
rect 119662 -6102 155426 -5866
rect 155662 -6102 191426 -5866
rect 191662 -6102 227426 -5866
rect 227662 -6102 263426 -5866
rect 263662 -6102 299426 -5866
rect 299662 -6102 335426 -5866
rect 335662 -6102 371426 -5866
rect 371662 -6102 407426 -5866
rect 407662 -6102 443426 -5866
rect 443662 -6102 479426 -5866
rect 479662 -6102 515426 -5866
rect 515662 -6102 551426 -5866
rect 551662 -6102 591022 -5866
rect 591258 -6102 591430 -5866
rect -7506 -6186 591430 -6102
rect -7506 -6422 -7334 -6186
rect -7098 -6422 11426 -6186
rect 11662 -6422 47426 -6186
rect 47662 -6422 83426 -6186
rect 83662 -6422 119426 -6186
rect 119662 -6422 155426 -6186
rect 155662 -6422 191426 -6186
rect 191662 -6422 227426 -6186
rect 227662 -6422 263426 -6186
rect 263662 -6422 299426 -6186
rect 299662 -6422 335426 -6186
rect 335662 -6422 371426 -6186
rect 371662 -6422 407426 -6186
rect 407662 -6422 443426 -6186
rect 443662 -6422 479426 -6186
rect 479662 -6422 515426 -6186
rect 515662 -6422 551426 -6186
rect 551662 -6422 591022 -6186
rect 591258 -6422 591430 -6186
rect -7506 -6434 591430 -6422
rect -7506 -6446 -6926 -6434
rect 11254 -6446 11834 -6434
rect 47254 -6446 47834 -6434
rect 83254 -6446 83834 -6434
rect 119254 -6446 119834 -6434
rect 155254 -6446 155834 -6434
rect 191254 -6446 191834 -6434
rect 227254 -6446 227834 -6434
rect 263254 -6446 263834 -6434
rect 299254 -6446 299834 -6434
rect 335254 -6446 335834 -6434
rect 371254 -6446 371834 -6434
rect 407254 -6446 407834 -6434
rect 443254 -6446 443834 -6434
rect 479254 -6446 479834 -6434
rect 515254 -6446 515834 -6434
rect 551254 -6446 551834 -6434
rect 590850 -6446 591430 -6434
rect -8426 -6774 -7846 -6762
rect 29254 -6774 29834 -6762
rect 65254 -6774 65834 -6762
rect 101254 -6774 101834 -6762
rect 137254 -6774 137834 -6762
rect 173254 -6774 173834 -6762
rect 209254 -6774 209834 -6762
rect 245254 -6774 245834 -6762
rect 281254 -6774 281834 -6762
rect 317254 -6774 317834 -6762
rect 353254 -6774 353834 -6762
rect 389254 -6774 389834 -6762
rect 425254 -6774 425834 -6762
rect 461254 -6774 461834 -6762
rect 497254 -6774 497834 -6762
rect 533254 -6774 533834 -6762
rect 569254 -6774 569834 -6762
rect 591770 -6774 592350 -6762
rect -8426 -6786 592350 -6774
rect -8426 -7022 -8254 -6786
rect -8018 -7022 29426 -6786
rect 29662 -7022 65426 -6786
rect 65662 -7022 101426 -6786
rect 101662 -7022 137426 -6786
rect 137662 -7022 173426 -6786
rect 173662 -7022 209426 -6786
rect 209662 -7022 245426 -6786
rect 245662 -7022 281426 -6786
rect 281662 -7022 317426 -6786
rect 317662 -7022 353426 -6786
rect 353662 -7022 389426 -6786
rect 389662 -7022 425426 -6786
rect 425662 -7022 461426 -6786
rect 461662 -7022 497426 -6786
rect 497662 -7022 533426 -6786
rect 533662 -7022 569426 -6786
rect 569662 -7022 591942 -6786
rect 592178 -7022 592350 -6786
rect -8426 -7106 592350 -7022
rect -8426 -7342 -8254 -7106
rect -8018 -7342 29426 -7106
rect 29662 -7342 65426 -7106
rect 65662 -7342 101426 -7106
rect 101662 -7342 137426 -7106
rect 137662 -7342 173426 -7106
rect 173662 -7342 209426 -7106
rect 209662 -7342 245426 -7106
rect 245662 -7342 281426 -7106
rect 281662 -7342 317426 -7106
rect 317662 -7342 353426 -7106
rect 353662 -7342 389426 -7106
rect 389662 -7342 425426 -7106
rect 425662 -7342 461426 -7106
rect 461662 -7342 497426 -7106
rect 497662 -7342 533426 -7106
rect 533662 -7342 569426 -7106
rect 569662 -7342 591942 -7106
rect 592178 -7342 592350 -7106
rect -8426 -7354 592350 -7342
rect -8426 -7366 -7846 -7354
rect 29254 -7366 29834 -7354
rect 65254 -7366 65834 -7354
rect 101254 -7366 101834 -7354
rect 137254 -7366 137834 -7354
rect 173254 -7366 173834 -7354
rect 209254 -7366 209834 -7354
rect 245254 -7366 245834 -7354
rect 281254 -7366 281834 -7354
rect 317254 -7366 317834 -7354
rect 353254 -7366 353834 -7354
rect 389254 -7366 389834 -7354
rect 425254 -7366 425834 -7354
rect 461254 -7366 461834 -7354
rect 497254 -7366 497834 -7354
rect 533254 -7366 533834 -7354
rect 569254 -7366 569834 -7354
rect 591770 -7366 592350 -7354
use rapcore  rapcore
timestamp 1607962800
transform 1 0 230200 0 1 340000
box 0 0 130000 130000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1986 -914 585910 -334 8 vccd1
port 636 nsew default input
rlabel metal5 s -2906 -1834 586830 -1254 8 vssd1
port 637 nsew default input
rlabel metal5 s -3826 -2754 587750 -2174 8 vccd2
port 638 nsew default input
rlabel metal5 s -4746 -3674 588670 -3094 8 vssd2
port 639 nsew default input
rlabel metal5 s -5666 -4594 589590 -4014 8 vdda1
port 640 nsew default input
rlabel metal5 s -6586 -5514 590510 -4934 8 vssa1
port 641 nsew default input
rlabel metal5 s -7506 -6434 591430 -5854 8 vdda2
port 642 nsew default input
rlabel metal5 s -8426 -7354 592350 -6774 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
