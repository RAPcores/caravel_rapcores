VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 2429.200 1573.130 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 1572.810 2429.060 2901.150 2429.200 ;
        RECT 1572.810 2429.000 1573.130 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 1568.210 2363.580 1568.530 2363.640 ;
        RECT 1572.810 2363.580 1573.130 2363.640 ;
        RECT 1568.210 2363.440 1573.130 2363.580 ;
        RECT 1568.210 2363.380 1568.530 2363.440 ;
        RECT 1572.810 2363.380 1573.130 2363.440 ;
      LAYER via ;
        RECT 1572.840 2429.000 1573.100 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 1568.240 2363.380 1568.500 2363.640 ;
        RECT 1572.840 2363.380 1573.100 2363.640 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 1572.840 2428.970 1573.100 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 1572.900 2363.670 1573.040 2428.970 ;
        RECT 1568.240 2363.350 1568.500 2363.670 ;
        RECT 1572.840 2363.350 1573.100 2363.670 ;
        RECT 1568.300 2350.000 1568.440 2363.350 ;
        RECT 1568.300 2349.740 1568.590 2350.000 ;
        RECT 1568.310 2346.000 1568.590 2349.740 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1821.745 2898.245 1821.915 2946.355 ;
        RECT 1822.205 2815.285 1822.375 2849.455 ;
      LAYER mcon ;
        RECT 1821.745 2946.185 1821.915 2946.355 ;
        RECT 1822.205 2849.285 1822.375 2849.455 ;
      LAYER met1 ;
        RECT 1821.670 3464.160 1821.990 3464.220 ;
        RECT 1825.350 3464.160 1825.670 3464.220 ;
        RECT 1821.670 3464.020 1825.670 3464.160 ;
        RECT 1821.670 3463.960 1821.990 3464.020 ;
        RECT 1825.350 3463.960 1825.670 3464.020 ;
        RECT 1821.670 3367.600 1821.990 3367.660 ;
        RECT 1822.590 3367.600 1822.910 3367.660 ;
        RECT 1821.670 3367.460 1822.910 3367.600 ;
        RECT 1821.670 3367.400 1821.990 3367.460 ;
        RECT 1822.590 3367.400 1822.910 3367.460 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1821.670 3174.140 1821.990 3174.200 ;
        RECT 1822.590 3174.140 1822.910 3174.200 ;
        RECT 1821.670 3174.000 1822.910 3174.140 ;
        RECT 1821.670 3173.940 1821.990 3174.000 ;
        RECT 1822.590 3173.940 1822.910 3174.000 ;
        RECT 1821.670 3077.580 1821.990 3077.640 ;
        RECT 1822.590 3077.580 1822.910 3077.640 ;
        RECT 1821.670 3077.440 1822.910 3077.580 ;
        RECT 1821.670 3077.380 1821.990 3077.440 ;
        RECT 1822.590 3077.380 1822.910 3077.440 ;
        RECT 1821.670 2981.020 1821.990 2981.080 ;
        RECT 1822.590 2981.020 1822.910 2981.080 ;
        RECT 1821.670 2980.880 1822.910 2981.020 ;
        RECT 1821.670 2980.820 1821.990 2980.880 ;
        RECT 1822.590 2980.820 1822.910 2980.880 ;
        RECT 1821.685 2946.340 1821.975 2946.385 ;
        RECT 1822.130 2946.340 1822.450 2946.400 ;
        RECT 1821.685 2946.200 1822.450 2946.340 ;
        RECT 1821.685 2946.155 1821.975 2946.200 ;
        RECT 1822.130 2946.140 1822.450 2946.200 ;
        RECT 1821.670 2898.400 1821.990 2898.460 ;
        RECT 1821.475 2898.260 1821.990 2898.400 ;
        RECT 1821.670 2898.200 1821.990 2898.260 ;
        RECT 1822.130 2849.440 1822.450 2849.500 ;
        RECT 1821.935 2849.300 1822.450 2849.440 ;
        RECT 1822.130 2849.240 1822.450 2849.300 ;
        RECT 1822.145 2815.440 1822.435 2815.485 ;
        RECT 1823.050 2815.440 1823.370 2815.500 ;
        RECT 1822.145 2815.300 1823.370 2815.440 ;
        RECT 1822.145 2815.255 1822.435 2815.300 ;
        RECT 1823.050 2815.240 1823.370 2815.300 ;
        RECT 1822.130 2753.220 1822.450 2753.280 ;
        RECT 1823.510 2753.220 1823.830 2753.280 ;
        RECT 1822.130 2753.080 1823.830 2753.220 ;
        RECT 1822.130 2753.020 1822.450 2753.080 ;
        RECT 1823.510 2753.020 1823.830 2753.080 ;
        RECT 1823.510 2719.220 1823.830 2719.280 ;
        RECT 1823.140 2719.080 1823.830 2719.220 ;
        RECT 1823.140 2718.600 1823.280 2719.080 ;
        RECT 1823.510 2719.020 1823.830 2719.080 ;
        RECT 1823.050 2718.340 1823.370 2718.600 ;
        RECT 1822.130 2656.660 1822.450 2656.720 ;
        RECT 1823.510 2656.660 1823.830 2656.720 ;
        RECT 1822.130 2656.520 1823.830 2656.660 ;
        RECT 1822.130 2656.460 1822.450 2656.520 ;
        RECT 1823.510 2656.460 1823.830 2656.520 ;
        RECT 1823.510 2622.660 1823.830 2622.720 ;
        RECT 1823.140 2622.520 1823.830 2622.660 ;
        RECT 1823.140 2622.040 1823.280 2622.520 ;
        RECT 1823.510 2622.460 1823.830 2622.520 ;
        RECT 1823.050 2621.780 1823.370 2622.040 ;
        RECT 1822.130 2560.100 1822.450 2560.160 ;
        RECT 1823.510 2560.100 1823.830 2560.160 ;
        RECT 1822.130 2559.960 1823.830 2560.100 ;
        RECT 1822.130 2559.900 1822.450 2559.960 ;
        RECT 1823.510 2559.900 1823.830 2559.960 ;
        RECT 1822.590 2511.820 1822.910 2511.880 ;
        RECT 1823.510 2511.820 1823.830 2511.880 ;
        RECT 1822.590 2511.680 1823.830 2511.820 ;
        RECT 1822.590 2511.620 1822.910 2511.680 ;
        RECT 1823.510 2511.620 1823.830 2511.680 ;
        RECT 1821.670 2401.320 1821.990 2401.380 ;
        RECT 1822.590 2401.320 1822.910 2401.380 ;
        RECT 1821.670 2401.180 1822.910 2401.320 ;
        RECT 1821.670 2401.120 1821.990 2401.180 ;
        RECT 1822.590 2401.120 1822.910 2401.180 ;
        RECT 1821.670 2304.760 1821.990 2304.820 ;
        RECT 1822.590 2304.760 1822.910 2304.820 ;
        RECT 1821.670 2304.620 1822.910 2304.760 ;
        RECT 1821.670 2304.560 1821.990 2304.620 ;
        RECT 1822.590 2304.560 1822.910 2304.620 ;
        RECT 1821.670 2208.200 1821.990 2208.260 ;
        RECT 1822.590 2208.200 1822.910 2208.260 ;
        RECT 1821.670 2208.060 1822.910 2208.200 ;
        RECT 1821.670 2208.000 1821.990 2208.060 ;
        RECT 1822.590 2208.000 1822.910 2208.060 ;
        RECT 1821.670 2111.640 1821.990 2111.700 ;
        RECT 1822.590 2111.640 1822.910 2111.700 ;
        RECT 1821.670 2111.500 1822.910 2111.640 ;
        RECT 1821.670 2111.440 1821.990 2111.500 ;
        RECT 1822.590 2111.440 1822.910 2111.500 ;
        RECT 1821.670 2015.080 1821.990 2015.140 ;
        RECT 1822.590 2015.080 1822.910 2015.140 ;
        RECT 1821.670 2014.940 1822.910 2015.080 ;
        RECT 1821.670 2014.880 1821.990 2014.940 ;
        RECT 1822.590 2014.880 1822.910 2014.940 ;
        RECT 1821.670 1918.520 1821.990 1918.580 ;
        RECT 1822.590 1918.520 1822.910 1918.580 ;
        RECT 1821.670 1918.380 1822.910 1918.520 ;
        RECT 1821.670 1918.320 1821.990 1918.380 ;
        RECT 1822.590 1918.320 1822.910 1918.380 ;
        RECT 1821.670 1821.960 1821.990 1822.020 ;
        RECT 1822.590 1821.960 1822.910 1822.020 ;
        RECT 1821.670 1821.820 1822.910 1821.960 ;
        RECT 1821.670 1821.760 1821.990 1821.820 ;
        RECT 1822.590 1821.760 1822.910 1821.820 ;
        RECT 1821.670 1725.400 1821.990 1725.460 ;
        RECT 1822.590 1725.400 1822.910 1725.460 ;
        RECT 1821.670 1725.260 1822.910 1725.400 ;
        RECT 1821.670 1725.200 1821.990 1725.260 ;
        RECT 1822.590 1725.200 1822.910 1725.260 ;
        RECT 1272.430 1689.360 1272.750 1689.420 ;
        RECT 1821.670 1689.360 1821.990 1689.420 ;
        RECT 1272.430 1689.220 1821.990 1689.360 ;
        RECT 1272.430 1689.160 1272.750 1689.220 ;
        RECT 1821.670 1689.160 1821.990 1689.220 ;
      LAYER via ;
        RECT 1821.700 3463.960 1821.960 3464.220 ;
        RECT 1825.380 3463.960 1825.640 3464.220 ;
        RECT 1821.700 3367.400 1821.960 3367.660 ;
        RECT 1822.620 3367.400 1822.880 3367.660 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1821.700 3173.940 1821.960 3174.200 ;
        RECT 1822.620 3173.940 1822.880 3174.200 ;
        RECT 1821.700 3077.380 1821.960 3077.640 ;
        RECT 1822.620 3077.380 1822.880 3077.640 ;
        RECT 1821.700 2980.820 1821.960 2981.080 ;
        RECT 1822.620 2980.820 1822.880 2981.080 ;
        RECT 1822.160 2946.140 1822.420 2946.400 ;
        RECT 1821.700 2898.200 1821.960 2898.460 ;
        RECT 1822.160 2849.240 1822.420 2849.500 ;
        RECT 1823.080 2815.240 1823.340 2815.500 ;
        RECT 1822.160 2753.020 1822.420 2753.280 ;
        RECT 1823.540 2753.020 1823.800 2753.280 ;
        RECT 1823.540 2719.020 1823.800 2719.280 ;
        RECT 1823.080 2718.340 1823.340 2718.600 ;
        RECT 1822.160 2656.460 1822.420 2656.720 ;
        RECT 1823.540 2656.460 1823.800 2656.720 ;
        RECT 1823.540 2622.460 1823.800 2622.720 ;
        RECT 1823.080 2621.780 1823.340 2622.040 ;
        RECT 1822.160 2559.900 1822.420 2560.160 ;
        RECT 1823.540 2559.900 1823.800 2560.160 ;
        RECT 1822.620 2511.620 1822.880 2511.880 ;
        RECT 1823.540 2511.620 1823.800 2511.880 ;
        RECT 1821.700 2401.120 1821.960 2401.380 ;
        RECT 1822.620 2401.120 1822.880 2401.380 ;
        RECT 1821.700 2304.560 1821.960 2304.820 ;
        RECT 1822.620 2304.560 1822.880 2304.820 ;
        RECT 1821.700 2208.000 1821.960 2208.260 ;
        RECT 1822.620 2208.000 1822.880 2208.260 ;
        RECT 1821.700 2111.440 1821.960 2111.700 ;
        RECT 1822.620 2111.440 1822.880 2111.700 ;
        RECT 1821.700 2014.880 1821.960 2015.140 ;
        RECT 1822.620 2014.880 1822.880 2015.140 ;
        RECT 1821.700 1918.320 1821.960 1918.580 ;
        RECT 1822.620 1918.320 1822.880 1918.580 ;
        RECT 1821.700 1821.760 1821.960 1822.020 ;
        RECT 1822.620 1821.760 1822.880 1822.020 ;
        RECT 1821.700 1725.200 1821.960 1725.460 ;
        RECT 1822.620 1725.200 1822.880 1725.460 ;
        RECT 1272.460 1689.160 1272.720 1689.420 ;
        RECT 1821.700 1689.160 1821.960 1689.420 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3464.250 1825.580 3517.230 ;
        RECT 1821.700 3463.930 1821.960 3464.250 ;
        RECT 1825.380 3463.930 1825.640 3464.250 ;
        RECT 1821.760 3415.370 1821.900 3463.930 ;
        RECT 1821.760 3415.230 1822.820 3415.370 ;
        RECT 1822.680 3367.690 1822.820 3415.230 ;
        RECT 1821.700 3367.370 1821.960 3367.690 ;
        RECT 1822.620 3367.370 1822.880 3367.690 ;
        RECT 1821.760 3318.810 1821.900 3367.370 ;
        RECT 1821.760 3318.670 1822.820 3318.810 ;
        RECT 1822.680 3270.790 1822.820 3318.670 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3222.250 1821.900 3270.470 ;
        RECT 1821.760 3222.110 1822.820 3222.250 ;
        RECT 1822.680 3174.230 1822.820 3222.110 ;
        RECT 1821.700 3173.910 1821.960 3174.230 ;
        RECT 1822.620 3173.910 1822.880 3174.230 ;
        RECT 1821.760 3125.690 1821.900 3173.910 ;
        RECT 1821.760 3125.550 1822.820 3125.690 ;
        RECT 1822.680 3077.670 1822.820 3125.550 ;
        RECT 1821.700 3077.350 1821.960 3077.670 ;
        RECT 1822.620 3077.350 1822.880 3077.670 ;
        RECT 1821.760 3029.130 1821.900 3077.350 ;
        RECT 1821.760 3028.990 1822.820 3029.130 ;
        RECT 1822.680 2981.110 1822.820 3028.990 ;
        RECT 1821.700 2980.850 1821.960 2981.110 ;
        RECT 1821.700 2980.790 1822.360 2980.850 ;
        RECT 1822.620 2980.790 1822.880 2981.110 ;
        RECT 1821.760 2980.710 1822.360 2980.790 ;
        RECT 1822.220 2980.170 1822.360 2980.710 ;
        RECT 1822.220 2980.030 1822.820 2980.170 ;
        RECT 1822.680 2959.770 1822.820 2980.030 ;
        RECT 1822.220 2959.630 1822.820 2959.770 ;
        RECT 1822.220 2946.430 1822.360 2959.630 ;
        RECT 1822.160 2946.110 1822.420 2946.430 ;
        RECT 1821.700 2898.170 1821.960 2898.490 ;
        RECT 1821.760 2863.210 1821.900 2898.170 ;
        RECT 1821.760 2863.070 1822.360 2863.210 ;
        RECT 1822.220 2849.530 1822.360 2863.070 ;
        RECT 1822.160 2849.210 1822.420 2849.530 ;
        RECT 1823.080 2815.210 1823.340 2815.530 ;
        RECT 1823.140 2801.445 1823.280 2815.210 ;
        RECT 1822.150 2801.075 1822.430 2801.445 ;
        RECT 1823.070 2801.075 1823.350 2801.445 ;
        RECT 1822.220 2753.310 1822.360 2801.075 ;
        RECT 1822.160 2752.990 1822.420 2753.310 ;
        RECT 1823.540 2752.990 1823.800 2753.310 ;
        RECT 1823.600 2719.310 1823.740 2752.990 ;
        RECT 1823.540 2718.990 1823.800 2719.310 ;
        RECT 1823.080 2718.310 1823.340 2718.630 ;
        RECT 1823.140 2704.885 1823.280 2718.310 ;
        RECT 1822.150 2704.515 1822.430 2704.885 ;
        RECT 1823.070 2704.515 1823.350 2704.885 ;
        RECT 1822.220 2656.750 1822.360 2704.515 ;
        RECT 1822.160 2656.430 1822.420 2656.750 ;
        RECT 1823.540 2656.430 1823.800 2656.750 ;
        RECT 1823.600 2622.750 1823.740 2656.430 ;
        RECT 1823.540 2622.430 1823.800 2622.750 ;
        RECT 1823.080 2621.750 1823.340 2622.070 ;
        RECT 1823.140 2608.325 1823.280 2621.750 ;
        RECT 1822.150 2607.955 1822.430 2608.325 ;
        RECT 1823.070 2607.955 1823.350 2608.325 ;
        RECT 1822.220 2560.190 1822.360 2607.955 ;
        RECT 1822.160 2559.870 1822.420 2560.190 ;
        RECT 1823.540 2559.870 1823.800 2560.190 ;
        RECT 1823.600 2511.910 1823.740 2559.870 ;
        RECT 1822.620 2511.765 1822.880 2511.910 ;
        RECT 1821.230 2511.395 1821.510 2511.765 ;
        RECT 1822.610 2511.395 1822.890 2511.765 ;
        RECT 1823.540 2511.590 1823.800 2511.910 ;
        RECT 1821.300 2463.485 1821.440 2511.395 ;
        RECT 1821.230 2463.115 1821.510 2463.485 ;
        RECT 1822.150 2463.115 1822.430 2463.485 ;
        RECT 1822.220 2449.770 1822.360 2463.115 ;
        RECT 1822.220 2449.630 1822.820 2449.770 ;
        RECT 1822.680 2401.410 1822.820 2449.630 ;
        RECT 1821.700 2401.090 1821.960 2401.410 ;
        RECT 1822.620 2401.090 1822.880 2401.410 ;
        RECT 1821.760 2400.810 1821.900 2401.090 ;
        RECT 1821.760 2400.670 1822.360 2400.810 ;
        RECT 1822.220 2353.210 1822.360 2400.670 ;
        RECT 1822.220 2353.070 1822.820 2353.210 ;
        RECT 1822.680 2304.850 1822.820 2353.070 ;
        RECT 1821.700 2304.530 1821.960 2304.850 ;
        RECT 1822.620 2304.530 1822.880 2304.850 ;
        RECT 1821.760 2304.250 1821.900 2304.530 ;
        RECT 1821.760 2304.110 1822.360 2304.250 ;
        RECT 1822.220 2256.650 1822.360 2304.110 ;
        RECT 1822.220 2256.510 1822.820 2256.650 ;
        RECT 1822.680 2208.290 1822.820 2256.510 ;
        RECT 1821.700 2207.970 1821.960 2208.290 ;
        RECT 1822.620 2207.970 1822.880 2208.290 ;
        RECT 1821.760 2207.690 1821.900 2207.970 ;
        RECT 1821.760 2207.550 1822.360 2207.690 ;
        RECT 1822.220 2160.090 1822.360 2207.550 ;
        RECT 1822.220 2159.950 1822.820 2160.090 ;
        RECT 1822.680 2111.730 1822.820 2159.950 ;
        RECT 1821.700 2111.410 1821.960 2111.730 ;
        RECT 1822.620 2111.410 1822.880 2111.730 ;
        RECT 1821.760 2111.130 1821.900 2111.410 ;
        RECT 1821.760 2110.990 1822.360 2111.130 ;
        RECT 1822.220 2063.530 1822.360 2110.990 ;
        RECT 1822.220 2063.390 1822.820 2063.530 ;
        RECT 1822.680 2015.170 1822.820 2063.390 ;
        RECT 1821.700 2014.850 1821.960 2015.170 ;
        RECT 1822.620 2014.850 1822.880 2015.170 ;
        RECT 1821.760 2014.570 1821.900 2014.850 ;
        RECT 1821.760 2014.430 1822.360 2014.570 ;
        RECT 1822.220 1966.970 1822.360 2014.430 ;
        RECT 1822.220 1966.830 1822.820 1966.970 ;
        RECT 1822.680 1918.610 1822.820 1966.830 ;
        RECT 1821.700 1918.290 1821.960 1918.610 ;
        RECT 1822.620 1918.290 1822.880 1918.610 ;
        RECT 1821.760 1918.010 1821.900 1918.290 ;
        RECT 1821.760 1917.870 1822.360 1918.010 ;
        RECT 1822.220 1870.410 1822.360 1917.870 ;
        RECT 1822.220 1870.270 1822.820 1870.410 ;
        RECT 1822.680 1822.050 1822.820 1870.270 ;
        RECT 1821.700 1821.730 1821.960 1822.050 ;
        RECT 1822.620 1821.730 1822.880 1822.050 ;
        RECT 1821.760 1773.170 1821.900 1821.730 ;
        RECT 1821.760 1773.030 1822.820 1773.170 ;
        RECT 1822.680 1725.490 1822.820 1773.030 ;
        RECT 1821.700 1725.170 1821.960 1725.490 ;
        RECT 1822.620 1725.170 1822.880 1725.490 ;
        RECT 1272.530 1700.340 1272.810 1704.000 ;
        RECT 1272.520 1700.000 1272.810 1700.340 ;
        RECT 1272.520 1689.450 1272.660 1700.000 ;
        RECT 1821.760 1689.450 1821.900 1725.170 ;
        RECT 1272.460 1689.130 1272.720 1689.450 ;
        RECT 1821.700 1689.130 1821.960 1689.450 ;
      LAYER via2 ;
        RECT 1822.150 2801.120 1822.430 2801.400 ;
        RECT 1823.070 2801.120 1823.350 2801.400 ;
        RECT 1822.150 2704.560 1822.430 2704.840 ;
        RECT 1823.070 2704.560 1823.350 2704.840 ;
        RECT 1822.150 2608.000 1822.430 2608.280 ;
        RECT 1823.070 2608.000 1823.350 2608.280 ;
        RECT 1821.230 2511.440 1821.510 2511.720 ;
        RECT 1822.610 2511.440 1822.890 2511.720 ;
        RECT 1821.230 2463.160 1821.510 2463.440 ;
        RECT 1822.150 2463.160 1822.430 2463.440 ;
      LAYER met3 ;
        RECT 1822.125 2801.410 1822.455 2801.425 ;
        RECT 1823.045 2801.410 1823.375 2801.425 ;
        RECT 1822.125 2801.110 1823.375 2801.410 ;
        RECT 1822.125 2801.095 1822.455 2801.110 ;
        RECT 1823.045 2801.095 1823.375 2801.110 ;
        RECT 1822.125 2704.850 1822.455 2704.865 ;
        RECT 1823.045 2704.850 1823.375 2704.865 ;
        RECT 1822.125 2704.550 1823.375 2704.850 ;
        RECT 1822.125 2704.535 1822.455 2704.550 ;
        RECT 1823.045 2704.535 1823.375 2704.550 ;
        RECT 1822.125 2608.290 1822.455 2608.305 ;
        RECT 1823.045 2608.290 1823.375 2608.305 ;
        RECT 1822.125 2607.990 1823.375 2608.290 ;
        RECT 1822.125 2607.975 1822.455 2607.990 ;
        RECT 1823.045 2607.975 1823.375 2607.990 ;
        RECT 1821.205 2511.730 1821.535 2511.745 ;
        RECT 1822.585 2511.730 1822.915 2511.745 ;
        RECT 1821.205 2511.430 1822.915 2511.730 ;
        RECT 1821.205 2511.415 1821.535 2511.430 ;
        RECT 1822.585 2511.415 1822.915 2511.430 ;
        RECT 1821.205 2463.450 1821.535 2463.465 ;
        RECT 1822.125 2463.450 1822.455 2463.465 ;
        RECT 1821.205 2463.150 1822.455 2463.450 ;
        RECT 1821.205 2463.135 1821.535 2463.150 ;
        RECT 1822.125 2463.135 1822.455 2463.150 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.010 3502.580 1145.330 3502.640 ;
        RECT 1500.590 3502.580 1500.910 3502.640 ;
        RECT 1145.010 3502.440 1500.910 3502.580 ;
        RECT 1145.010 3502.380 1145.330 3502.440 ;
        RECT 1500.590 3502.380 1500.910 3502.440 ;
      LAYER via ;
        RECT 1145.040 3502.380 1145.300 3502.640 ;
        RECT 1500.620 3502.380 1500.880 3502.640 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3502.670 1500.820 3517.600 ;
        RECT 1145.040 3502.350 1145.300 3502.670 ;
        RECT 1500.620 3502.350 1500.880 3502.670 ;
        RECT 1145.100 2024.885 1145.240 3502.350 ;
        RECT 1145.030 2024.515 1145.310 2024.885 ;
      LAYER via2 ;
        RECT 1145.030 2024.560 1145.310 2024.840 ;
      LAYER met3 ;
        RECT 1145.005 2024.850 1145.335 2024.865 ;
        RECT 1151.000 2024.850 1155.000 2025.000 ;
        RECT 1145.005 2024.550 1155.000 2024.850 ;
        RECT 1145.005 2024.535 1145.335 2024.550 ;
        RECT 1151.000 2024.400 1155.000 2024.550 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 1690.380 17.870 1690.440 ;
        RECT 1760.030 1690.380 1760.350 1690.440 ;
        RECT 17.550 1690.240 1760.350 1690.380 ;
        RECT 17.550 1690.180 17.870 1690.240 ;
        RECT 1760.030 1690.180 1760.350 1690.240 ;
      LAYER via ;
        RECT 17.580 1690.180 17.840 1690.440 ;
        RECT 1760.060 1690.180 1760.320 1690.440 ;
      LAYER met2 ;
        RECT 17.570 3124.075 17.850 3124.445 ;
        RECT 17.640 1690.470 17.780 3124.075 ;
        RECT 1760.130 1700.340 1760.410 1704.000 ;
        RECT 1760.120 1700.000 1760.410 1700.340 ;
        RECT 1760.120 1690.470 1760.260 1700.000 ;
        RECT 17.580 1690.150 17.840 1690.470 ;
        RECT 1760.060 1690.150 1760.320 1690.470 ;
      LAYER via2 ;
        RECT 17.570 3124.120 17.850 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.545 3124.410 17.875 3124.425 ;
        RECT -4.800 3124.110 17.875 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.545 3124.095 17.875 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2836.180 16.950 2836.240 ;
        RECT 1794.990 2836.180 1795.310 2836.240 ;
        RECT 16.630 2836.040 1795.310 2836.180 ;
        RECT 16.630 2835.980 16.950 2836.040 ;
        RECT 1794.990 2835.980 1795.310 2836.040 ;
      LAYER via ;
        RECT 16.660 2835.980 16.920 2836.240 ;
        RECT 1795.020 2835.980 1795.280 2836.240 ;
      LAYER met2 ;
        RECT 16.650 2836.435 16.930 2836.805 ;
        RECT 16.720 2836.270 16.860 2836.435 ;
        RECT 16.660 2835.950 16.920 2836.270 ;
        RECT 1795.020 2835.950 1795.280 2836.270 ;
        RECT 1795.080 2243.730 1795.220 2835.950 ;
        RECT 1797.770 2243.730 1798.050 2243.845 ;
        RECT 1795.080 2243.590 1798.050 2243.730 ;
        RECT 1797.770 2243.475 1798.050 2243.590 ;
      LAYER via2 ;
        RECT 16.650 2836.480 16.930 2836.760 ;
        RECT 1797.770 2243.520 1798.050 2243.800 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 16.625 2836.770 16.955 2836.785 ;
        RECT -4.800 2836.470 16.955 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 16.625 2836.455 16.955 2836.470 ;
        RECT 1797.745 2243.810 1798.075 2243.825 ;
        RECT 1797.745 2243.495 1798.290 2243.810 ;
        RECT 1797.990 2241.920 1798.290 2243.495 ;
        RECT 1797.000 2241.320 1801.000 2241.920 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 1980.060 16.950 1980.120 ;
        RECT 1141.790 1980.060 1142.110 1980.120 ;
        RECT 16.630 1979.920 1086.820 1980.060 ;
        RECT 16.630 1979.860 16.950 1979.920 ;
        RECT 1086.680 1979.720 1086.820 1979.920 ;
        RECT 1094.960 1979.920 1142.110 1980.060 ;
        RECT 1094.960 1979.720 1095.100 1979.920 ;
        RECT 1141.790 1979.860 1142.110 1979.920 ;
        RECT 1086.680 1979.580 1095.100 1979.720 ;
      LAYER via ;
        RECT 16.660 1979.860 16.920 1980.120 ;
        RECT 1141.820 1979.860 1142.080 1980.120 ;
      LAYER met2 ;
        RECT 1141.810 2241.435 1142.090 2241.805 ;
        RECT 1141.880 1980.150 1142.020 2241.435 ;
        RECT 16.660 1979.830 16.920 1980.150 ;
        RECT 1141.820 1979.830 1142.080 1980.150 ;
        RECT 16.720 1975.245 16.860 1979.830 ;
        RECT 16.650 1974.875 16.930 1975.245 ;
      LAYER via2 ;
        RECT 1141.810 2241.480 1142.090 2241.760 ;
        RECT 16.650 1974.920 16.930 1975.200 ;
      LAYER met3 ;
        RECT 1141.785 2241.770 1142.115 2241.785 ;
        RECT 1151.000 2241.770 1155.000 2241.920 ;
        RECT 1141.785 2241.470 1155.000 2241.770 ;
        RECT 1141.785 2241.455 1142.115 2241.470 ;
        RECT 1151.000 2241.320 1155.000 2241.470 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 16.625 1975.210 16.955 1975.225 ;
        RECT -4.800 1974.910 16.955 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 16.625 1974.895 16.955 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.150 2359.755 1661.430 2360.125 ;
        RECT 1661.220 2350.000 1661.360 2359.755 ;
        RECT 1661.220 2349.740 1661.510 2350.000 ;
        RECT 1661.230 2346.000 1661.510 2349.740 ;
        RECT 17.110 1262.235 17.390 1262.605 ;
        RECT 17.180 1256.485 17.320 1262.235 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
      LAYER via2 ;
        RECT 1661.150 2359.800 1661.430 2360.080 ;
        RECT 17.110 1262.280 17.390 1262.560 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
      LAYER met3 ;
        RECT 1341.630 2360.090 1342.010 2360.100 ;
        RECT 1661.125 2360.090 1661.455 2360.105 ;
        RECT 1341.630 2359.790 1661.455 2360.090 ;
        RECT 1341.630 2359.780 1342.010 2359.790 ;
        RECT 1661.125 2359.775 1661.455 2359.790 ;
        RECT 17.085 1262.570 17.415 1262.585 ;
        RECT 1341.630 1262.570 1342.010 1262.580 ;
        RECT 17.085 1262.270 1342.010 1262.570 ;
        RECT 17.085 1262.255 17.415 1262.270 ;
        RECT 1341.630 1262.260 1342.010 1262.270 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
      LAYER via3 ;
        RECT 1341.660 2359.780 1341.980 2360.100 ;
        RECT 1341.660 1262.260 1341.980 1262.580 ;
      LAYER met4 ;
        RECT 1341.655 2359.775 1341.985 2360.105 ;
        RECT 1341.670 1262.585 1341.970 2359.775 ;
        RECT 1341.655 1262.255 1341.985 1262.585 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 2360.520 18.330 2360.580 ;
        RECT 1289.450 2360.520 1289.770 2360.580 ;
        RECT 18.010 2360.380 1289.770 2360.520 ;
        RECT 18.010 2360.320 18.330 2360.380 ;
        RECT 1289.450 2360.320 1289.770 2360.380 ;
      LAYER via ;
        RECT 18.040 2360.320 18.300 2360.580 ;
        RECT 1289.480 2360.320 1289.740 2360.580 ;
      LAYER met2 ;
        RECT 18.040 2360.290 18.300 2360.610 ;
        RECT 1289.480 2360.290 1289.740 2360.610 ;
        RECT 18.100 1040.925 18.240 2360.290 ;
        RECT 1289.540 2350.000 1289.680 2360.290 ;
        RECT 1289.540 2349.740 1289.830 2350.000 ;
        RECT 1289.550 2346.000 1289.830 2349.740 ;
        RECT 18.030 1040.555 18.310 1040.925 ;
      LAYER via2 ;
        RECT 18.030 1040.600 18.310 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 18.005 1040.890 18.335 1040.905 ;
        RECT -4.800 1040.590 18.335 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 18.005 1040.575 18.335 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2901.310 1964.675 2901.590 1965.045 ;
        RECT 2901.380 1814.765 2901.520 1964.675 ;
        RECT 2901.310 1814.395 2901.590 1814.765 ;
      LAYER via2 ;
        RECT 2901.310 1964.720 2901.590 1965.000 ;
        RECT 2901.310 1814.440 2901.590 1814.720 ;
      LAYER met3 ;
        RECT 2901.285 1965.010 2901.615 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2901.285 1964.710 2924.800 1965.010 ;
        RECT 2901.285 1964.695 2901.615 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 1797.950 1814.730 1798.330 1814.740 ;
        RECT 2901.285 1814.730 2901.615 1814.745 ;
        RECT 1797.950 1814.430 2901.615 1814.730 ;
        RECT 1797.950 1814.420 1798.330 1814.430 ;
        RECT 2901.285 1814.415 2901.615 1814.430 ;
        RECT 1151.000 1808.160 1155.000 1808.760 ;
        RECT 1153.990 1805.900 1154.290 1808.160 ;
        RECT 1153.950 1805.580 1154.330 1805.900 ;
      LAYER via3 ;
        RECT 1797.980 1814.420 1798.300 1814.740 ;
        RECT 1153.980 1805.580 1154.300 1805.900 ;
      LAYER met4 ;
        RECT 1194.950 1816.710 1196.130 1817.890 ;
        RECT 1242.790 1816.710 1243.970 1817.890 ;
        RECT 1343.990 1816.710 1345.170 1817.890 ;
        RECT 1723.950 1816.710 1725.130 1817.890 ;
        RECT 1153.975 1805.575 1154.305 1805.905 ;
        RECT 1153.990 1804.290 1154.290 1805.575 ;
        RECT 1195.390 1804.290 1195.690 1816.710 ;
        RECT 1243.230 1804.290 1243.530 1816.710 ;
        RECT 1344.430 1804.290 1344.730 1816.710 ;
        RECT 1724.390 1804.290 1724.690 1816.710 ;
        RECT 1797.975 1814.415 1798.305 1814.745 ;
        RECT 1797.990 1804.290 1798.290 1814.415 ;
        RECT 1153.550 1803.110 1154.730 1804.290 ;
        RECT 1194.950 1803.110 1196.130 1804.290 ;
        RECT 1242.790 1803.110 1243.970 1804.290 ;
        RECT 1343.990 1803.110 1345.170 1804.290 ;
        RECT 1723.950 1803.110 1725.130 1804.290 ;
        RECT 1797.550 1803.110 1798.730 1804.290 ;
      LAYER met5 ;
        RECT 1194.740 1816.500 1244.180 1818.100 ;
        RECT 1343.780 1816.500 1725.340 1818.100 ;
        RECT 1153.340 1802.900 1196.340 1804.500 ;
        RECT 1242.580 1802.900 1345.380 1804.500 ;
        RECT 1723.740 1802.900 1798.940 1804.500 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1797.290 2194.600 1797.610 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 1797.290 2194.460 2901.150 2194.600 ;
        RECT 1797.290 2194.400 1797.610 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
        RECT 1191.470 1689.700 1191.790 1689.760 ;
        RECT 1797.290 1689.700 1797.610 1689.760 ;
        RECT 1191.470 1689.560 1797.610 1689.700 ;
        RECT 1191.470 1689.500 1191.790 1689.560 ;
        RECT 1797.290 1689.500 1797.610 1689.560 ;
      LAYER via ;
        RECT 1797.320 2194.400 1797.580 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
        RECT 1191.500 1689.500 1191.760 1689.760 ;
        RECT 1797.320 1689.500 1797.580 1689.760 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 1797.320 2194.370 1797.580 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 1191.570 1700.340 1191.850 1704.000 ;
        RECT 1191.560 1700.000 1191.850 1700.340 ;
        RECT 1191.560 1689.790 1191.700 1700.000 ;
        RECT 1797.380 1689.790 1797.520 2194.370 ;
        RECT 1191.500 1689.470 1191.760 1689.790 ;
        RECT 1797.320 1689.470 1797.580 1689.790 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1812.010 2725.680 1812.330 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 1812.010 2725.540 2901.150 2725.680 ;
        RECT 1812.010 2725.480 1812.330 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 1812.040 2725.480 1812.300 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 1812.040 2725.450 1812.300 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 1812.100 1808.645 1812.240 2725.450 ;
        RECT 1812.030 1808.275 1812.310 1808.645 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 1812.030 1808.320 1812.310 1808.600 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 1797.000 1808.610 1801.000 1808.760 ;
        RECT 1812.005 1808.610 1812.335 1808.625 ;
        RECT 1797.000 1808.310 1812.335 1808.610 ;
        RECT 1797.000 1808.160 1801.000 1808.310 ;
        RECT 1812.005 1808.295 1812.335 1808.310 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1811.550 2960.280 1811.870 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1811.550 2960.140 2901.150 2960.280 ;
        RECT 1811.550 2960.080 1811.870 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 1811.580 2960.080 1811.840 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1811.580 2960.050 1811.840 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1811.640 1736.565 1811.780 2960.050 ;
        RECT 1811.570 1736.195 1811.850 1736.565 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 1811.570 1736.240 1811.850 1736.520 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 1797.000 1736.530 1801.000 1736.680 ;
        RECT 1811.545 1736.530 1811.875 1736.545 ;
        RECT 1797.000 1736.230 1811.875 1736.530 ;
        RECT 1797.000 1736.080 1801.000 1736.230 ;
        RECT 1811.545 1736.215 1811.875 1736.230 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1811.090 3429.480 1811.410 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 1811.090 3429.340 2901.150 3429.480 ;
        RECT 1811.090 3429.280 1811.410 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1811.120 3429.280 1811.380 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1811.120 3429.250 1811.380 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1811.180 2169.725 1811.320 3429.250 ;
        RECT 1811.110 2169.355 1811.390 2169.725 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 1811.110 2169.400 1811.390 2169.680 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 1797.000 2169.690 1801.000 2169.840 ;
        RECT 1811.085 2169.690 1811.415 2169.705 ;
        RECT 1797.000 2169.390 1811.415 2169.690 ;
        RECT 1797.000 2169.240 1801.000 2169.390 ;
        RECT 1811.085 2169.375 1811.415 2169.390 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1200.210 3501.900 1200.530 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 1200.210 3501.760 2717.610 3501.900 ;
        RECT 1200.210 3501.700 1200.530 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 1200.240 3501.700 1200.500 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 1200.240 3501.670 1200.500 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 1200.300 2350.490 1200.440 3501.670 ;
        RECT 1199.380 2350.350 1200.440 2350.490 ;
        RECT 1197.090 2349.130 1197.370 2350.000 ;
        RECT 1199.380 2349.130 1199.520 2350.350 ;
        RECT 1197.090 2348.990 1199.520 2349.130 ;
        RECT 1197.090 2346.000 1197.370 2348.990 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1817.990 3501.560 1818.310 3501.620 ;
        RECT 2392.530 3501.560 2392.850 3501.620 ;
        RECT 1817.990 3501.420 2392.850 3501.560 ;
        RECT 1817.990 3501.360 1818.310 3501.420 ;
        RECT 2392.530 3501.360 2392.850 3501.420 ;
        RECT 1434.810 1690.040 1435.130 1690.100 ;
        RECT 1817.990 1690.040 1818.310 1690.100 ;
        RECT 1434.810 1689.900 1818.310 1690.040 ;
        RECT 1434.810 1689.840 1435.130 1689.900 ;
        RECT 1817.990 1689.840 1818.310 1689.900 ;
      LAYER via ;
        RECT 1818.020 3501.360 1818.280 3501.620 ;
        RECT 2392.560 3501.360 2392.820 3501.620 ;
        RECT 1434.840 1689.840 1435.100 1690.100 ;
        RECT 1818.020 1689.840 1818.280 1690.100 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.650 2392.760 3517.600 ;
        RECT 1818.020 3501.330 1818.280 3501.650 ;
        RECT 2392.560 3501.330 2392.820 3501.650 ;
        RECT 1434.910 1700.340 1435.190 1704.000 ;
        RECT 1434.900 1700.000 1435.190 1700.340 ;
        RECT 1434.900 1690.130 1435.040 1700.000 ;
        RECT 1818.080 1690.130 1818.220 3501.330 ;
        RECT 1434.840 1689.810 1435.100 1690.130 ;
        RECT 1818.020 1689.810 1818.280 1690.130 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1831.790 3502.240 1832.110 3502.300 ;
        RECT 2068.230 3502.240 2068.550 3502.300 ;
        RECT 1831.790 3502.100 2068.550 3502.240 ;
        RECT 1831.790 3502.040 1832.110 3502.100 ;
        RECT 2068.230 3502.040 2068.550 3502.100 ;
        RECT 1597.650 1689.020 1597.970 1689.080 ;
        RECT 1831.790 1689.020 1832.110 1689.080 ;
        RECT 1597.650 1688.880 1832.110 1689.020 ;
        RECT 1597.650 1688.820 1597.970 1688.880 ;
        RECT 1831.790 1688.820 1832.110 1688.880 ;
      LAYER via ;
        RECT 1831.820 3502.040 1832.080 3502.300 ;
        RECT 2068.260 3502.040 2068.520 3502.300 ;
        RECT 1597.680 1688.820 1597.940 1689.080 ;
        RECT 1831.820 1688.820 1832.080 1689.080 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3502.330 2068.460 3517.600 ;
        RECT 1831.820 3502.010 1832.080 3502.330 ;
        RECT 2068.260 3502.010 2068.520 3502.330 ;
        RECT 1597.750 1700.340 1598.030 1704.000 ;
        RECT 1597.740 1700.000 1598.030 1700.340 ;
        RECT 1597.740 1689.110 1597.880 1700.000 ;
        RECT 1831.880 1689.110 1832.020 3502.010 ;
        RECT 1597.680 1688.790 1597.940 1689.110 ;
        RECT 1831.820 1688.790 1832.080 1689.110 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1476.210 3502.920 1476.530 3502.980 ;
        RECT 1743.930 3502.920 1744.250 3502.980 ;
        RECT 1476.210 3502.780 1744.250 3502.920 ;
        RECT 1476.210 3502.720 1476.530 3502.780 ;
        RECT 1743.930 3502.720 1744.250 3502.780 ;
      LAYER via ;
        RECT 1476.240 3502.720 1476.500 3502.980 ;
        RECT 1743.960 3502.720 1744.220 3502.980 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3503.010 1744.160 3517.600 ;
        RECT 1476.240 3502.690 1476.500 3503.010 ;
        RECT 1743.960 3502.690 1744.220 3503.010 ;
        RECT 1475.390 2349.810 1475.670 2350.000 ;
        RECT 1476.300 2349.810 1476.440 3502.690 ;
        RECT 1475.390 2349.670 1476.440 2349.810 ;
        RECT 1475.390 2346.000 1475.670 2349.670 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3502.240 1419.490 3502.300 ;
        RECT 1794.530 3502.240 1794.850 3502.300 ;
        RECT 1419.170 3502.100 1794.850 3502.240 ;
        RECT 1419.170 3502.040 1419.490 3502.100 ;
        RECT 1794.530 3502.040 1794.850 3502.100 ;
        RECT 1795.910 2096.680 1796.230 2096.740 ;
        RECT 1797.750 2096.680 1798.070 2096.740 ;
        RECT 1795.910 2096.540 1798.070 2096.680 ;
        RECT 1795.910 2096.480 1796.230 2096.540 ;
        RECT 1797.750 2096.480 1798.070 2096.540 ;
      LAYER via ;
        RECT 1419.200 3502.040 1419.460 3502.300 ;
        RECT 1794.560 3502.040 1794.820 3502.300 ;
        RECT 1795.940 2096.480 1796.200 2096.740 ;
        RECT 1797.780 2096.480 1798.040 2096.740 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3502.330 1419.400 3517.600 ;
        RECT 1419.200 3502.010 1419.460 3502.330 ;
        RECT 1794.560 3502.010 1794.820 3502.330 ;
        RECT 1794.620 2096.850 1794.760 3502.010 ;
        RECT 1794.620 2096.770 1796.140 2096.850 ;
        RECT 1794.620 2096.710 1796.200 2096.770 ;
        RECT 1795.940 2096.450 1796.200 2096.710 ;
        RECT 1797.780 2096.450 1798.040 2096.770 ;
        RECT 1797.840 2096.285 1797.980 2096.450 ;
        RECT 1797.770 2095.915 1798.050 2096.285 ;
      LAYER via2 ;
        RECT 1797.770 2095.960 1798.050 2096.240 ;
      LAYER met3 ;
        RECT 1797.000 2097.160 1801.000 2097.760 ;
        RECT 1797.990 2096.265 1798.290 2097.160 ;
        RECT 1797.745 2095.950 1798.290 2096.265 ;
        RECT 1797.745 2095.935 1798.075 2095.950 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1094.945 3332.765 1095.115 3380.875 ;
        RECT 1096.325 3236.205 1096.495 3284.315 ;
        RECT 1096.785 3084.225 1096.955 3132.675 ;
        RECT 1095.405 3043.425 1095.575 3057.195 ;
        RECT 1096.325 3007.725 1096.495 3042.915 ;
        RECT 1095.865 2946.525 1096.035 2994.635 ;
        RECT 1094.485 2849.625 1094.655 2898.075 ;
        RECT 1094.485 2753.065 1094.655 2767.175 ;
        RECT 1094.485 1980.245 1094.655 2028.355 ;
        RECT 1094.025 1773.865 1094.195 1801.235 ;
        RECT 1094.945 1752.105 1095.115 1773.355 ;
      LAYER mcon ;
        RECT 1094.945 3380.705 1095.115 3380.875 ;
        RECT 1096.325 3284.145 1096.495 3284.315 ;
        RECT 1096.785 3132.505 1096.955 3132.675 ;
        RECT 1095.405 3057.025 1095.575 3057.195 ;
        RECT 1096.325 3042.745 1096.495 3042.915 ;
        RECT 1095.865 2994.465 1096.035 2994.635 ;
        RECT 1094.485 2897.905 1094.655 2898.075 ;
        RECT 1094.485 2767.005 1094.655 2767.175 ;
        RECT 1094.485 2028.185 1094.655 2028.355 ;
        RECT 1094.025 1801.065 1094.195 1801.235 ;
        RECT 1094.945 1773.185 1095.115 1773.355 ;
      LAYER met1 ;
        RECT 1094.870 3470.960 1095.190 3471.020 ;
        RECT 1095.790 3470.960 1096.110 3471.020 ;
        RECT 1094.870 3470.820 1096.110 3470.960 ;
        RECT 1094.870 3470.760 1095.190 3470.820 ;
        RECT 1095.790 3470.760 1096.110 3470.820 ;
        RECT 1095.790 3443.420 1096.110 3443.480 ;
        RECT 1095.420 3443.280 1096.110 3443.420 ;
        RECT 1095.420 3443.140 1095.560 3443.280 ;
        RECT 1095.790 3443.220 1096.110 3443.280 ;
        RECT 1095.330 3442.880 1095.650 3443.140 ;
        RECT 1094.870 3380.860 1095.190 3380.920 ;
        RECT 1094.675 3380.720 1095.190 3380.860 ;
        RECT 1094.870 3380.660 1095.190 3380.720 ;
        RECT 1094.885 3332.920 1095.175 3332.965 ;
        RECT 1095.330 3332.920 1095.650 3332.980 ;
        RECT 1094.885 3332.780 1095.650 3332.920 ;
        RECT 1094.885 3332.735 1095.175 3332.780 ;
        RECT 1095.330 3332.720 1095.650 3332.780 ;
        RECT 1095.790 3298.240 1096.110 3298.300 ;
        RECT 1096.710 3298.240 1097.030 3298.300 ;
        RECT 1095.790 3298.100 1097.030 3298.240 ;
        RECT 1095.790 3298.040 1096.110 3298.100 ;
        RECT 1096.710 3298.040 1097.030 3298.100 ;
        RECT 1096.265 3284.300 1096.555 3284.345 ;
        RECT 1096.710 3284.300 1097.030 3284.360 ;
        RECT 1096.265 3284.160 1097.030 3284.300 ;
        RECT 1096.265 3284.115 1096.555 3284.160 ;
        RECT 1096.710 3284.100 1097.030 3284.160 ;
        RECT 1096.250 3236.360 1096.570 3236.420 ;
        RECT 1096.055 3236.220 1096.570 3236.360 ;
        RECT 1096.250 3236.160 1096.570 3236.220 ;
        RECT 1096.250 3202.020 1096.570 3202.080 ;
        RECT 1095.420 3201.880 1096.570 3202.020 ;
        RECT 1095.420 3201.400 1095.560 3201.880 ;
        RECT 1096.250 3201.820 1096.570 3201.880 ;
        RECT 1095.330 3201.140 1095.650 3201.400 ;
        RECT 1095.330 3187.740 1095.650 3187.800 ;
        RECT 1095.790 3187.740 1096.110 3187.800 ;
        RECT 1095.330 3187.600 1096.110 3187.740 ;
        RECT 1095.330 3187.540 1095.650 3187.600 ;
        RECT 1095.790 3187.540 1096.110 3187.600 ;
        RECT 1096.710 3132.660 1097.030 3132.720 ;
        RECT 1096.515 3132.520 1097.030 3132.660 ;
        RECT 1096.710 3132.460 1097.030 3132.520 ;
        RECT 1096.710 3084.380 1097.030 3084.440 ;
        RECT 1096.515 3084.240 1097.030 3084.380 ;
        RECT 1096.710 3084.180 1097.030 3084.240 ;
        RECT 1095.345 3057.180 1095.635 3057.225 ;
        RECT 1096.710 3057.180 1097.030 3057.240 ;
        RECT 1095.345 3057.040 1097.030 3057.180 ;
        RECT 1095.345 3056.995 1095.635 3057.040 ;
        RECT 1096.710 3056.980 1097.030 3057.040 ;
        RECT 1095.330 3043.580 1095.650 3043.640 ;
        RECT 1095.135 3043.440 1095.650 3043.580 ;
        RECT 1095.330 3043.380 1095.650 3043.440 ;
        RECT 1095.330 3042.900 1095.650 3042.960 ;
        RECT 1096.265 3042.900 1096.555 3042.945 ;
        RECT 1095.330 3042.760 1096.555 3042.900 ;
        RECT 1095.330 3042.700 1095.650 3042.760 ;
        RECT 1096.265 3042.715 1096.555 3042.760 ;
        RECT 1096.250 3007.880 1096.570 3007.940 ;
        RECT 1096.055 3007.740 1096.570 3007.880 ;
        RECT 1096.250 3007.680 1096.570 3007.740 ;
        RECT 1095.805 2994.620 1096.095 2994.665 ;
        RECT 1096.250 2994.620 1096.570 2994.680 ;
        RECT 1095.805 2994.480 1096.570 2994.620 ;
        RECT 1095.805 2994.435 1096.095 2994.480 ;
        RECT 1096.250 2994.420 1096.570 2994.480 ;
        RECT 1095.790 2946.680 1096.110 2946.740 ;
        RECT 1095.595 2946.540 1096.110 2946.680 ;
        RECT 1095.790 2946.480 1096.110 2946.540 ;
        RECT 1094.870 2912.000 1095.190 2912.060 ;
        RECT 1095.790 2912.000 1096.110 2912.060 ;
        RECT 1094.870 2911.860 1096.110 2912.000 ;
        RECT 1094.870 2911.800 1095.190 2911.860 ;
        RECT 1095.790 2911.800 1096.110 2911.860 ;
        RECT 1094.425 2898.060 1094.715 2898.105 ;
        RECT 1094.870 2898.060 1095.190 2898.120 ;
        RECT 1094.425 2897.920 1095.190 2898.060 ;
        RECT 1094.425 2897.875 1094.715 2897.920 ;
        RECT 1094.870 2897.860 1095.190 2897.920 ;
        RECT 1094.410 2849.780 1094.730 2849.840 ;
        RECT 1094.215 2849.640 1094.730 2849.780 ;
        RECT 1094.410 2849.580 1094.730 2849.640 ;
        RECT 1094.410 2815.240 1094.730 2815.500 ;
        RECT 1094.500 2814.760 1094.640 2815.240 ;
        RECT 1094.870 2814.760 1095.190 2814.820 ;
        RECT 1094.500 2814.620 1095.190 2814.760 ;
        RECT 1094.870 2814.560 1095.190 2814.620 ;
        RECT 1094.410 2767.160 1094.730 2767.220 ;
        RECT 1094.215 2767.020 1094.730 2767.160 ;
        RECT 1094.410 2766.960 1094.730 2767.020 ;
        RECT 1094.410 2753.220 1094.730 2753.280 ;
        RECT 1094.215 2753.080 1094.730 2753.220 ;
        RECT 1094.410 2753.020 1094.730 2753.080 ;
        RECT 1094.410 2718.680 1094.730 2718.940 ;
        RECT 1094.500 2718.200 1094.640 2718.680 ;
        RECT 1094.870 2718.200 1095.190 2718.260 ;
        RECT 1094.500 2718.060 1095.190 2718.200 ;
        RECT 1094.870 2718.000 1095.190 2718.060 ;
        RECT 1094.870 2621.640 1095.190 2621.700 ;
        RECT 1095.790 2621.640 1096.110 2621.700 ;
        RECT 1094.870 2621.500 1096.110 2621.640 ;
        RECT 1094.870 2621.440 1095.190 2621.500 ;
        RECT 1095.790 2621.440 1096.110 2621.500 ;
        RECT 1094.410 2511.820 1094.730 2511.880 ;
        RECT 1096.710 2511.820 1097.030 2511.880 ;
        RECT 1094.410 2511.680 1097.030 2511.820 ;
        RECT 1094.410 2511.620 1094.730 2511.680 ;
        RECT 1096.710 2511.620 1097.030 2511.680 ;
        RECT 1095.790 2401.320 1096.110 2401.380 ;
        RECT 1096.710 2401.320 1097.030 2401.380 ;
        RECT 1095.790 2401.180 1097.030 2401.320 ;
        RECT 1095.790 2401.120 1096.110 2401.180 ;
        RECT 1096.710 2401.120 1097.030 2401.180 ;
        RECT 1095.790 2304.760 1096.110 2304.820 ;
        RECT 1096.710 2304.760 1097.030 2304.820 ;
        RECT 1095.790 2304.620 1097.030 2304.760 ;
        RECT 1095.790 2304.560 1096.110 2304.620 ;
        RECT 1096.710 2304.560 1097.030 2304.620 ;
        RECT 1096.250 2221.800 1096.570 2221.860 ;
        RECT 1097.170 2221.800 1097.490 2221.860 ;
        RECT 1096.250 2221.660 1097.490 2221.800 ;
        RECT 1096.250 2221.600 1096.570 2221.660 ;
        RECT 1097.170 2221.600 1097.490 2221.660 ;
        RECT 1094.870 2139.180 1095.190 2139.240 ;
        RECT 1095.790 2139.180 1096.110 2139.240 ;
        RECT 1094.870 2139.040 1096.110 2139.180 ;
        RECT 1094.870 2138.980 1095.190 2139.040 ;
        RECT 1095.790 2138.980 1096.110 2139.040 ;
        RECT 1093.490 2125.240 1093.810 2125.300 ;
        RECT 1094.870 2125.240 1095.190 2125.300 ;
        RECT 1093.490 2125.100 1095.190 2125.240 ;
        RECT 1093.490 2125.040 1093.810 2125.100 ;
        RECT 1094.870 2125.040 1095.190 2125.100 ;
        RECT 1094.410 2042.420 1094.730 2042.680 ;
        RECT 1094.500 2041.940 1094.640 2042.420 ;
        RECT 1094.870 2041.940 1095.190 2042.000 ;
        RECT 1094.500 2041.800 1095.190 2041.940 ;
        RECT 1094.870 2041.740 1095.190 2041.800 ;
        RECT 1094.425 2028.340 1094.715 2028.385 ;
        RECT 1094.870 2028.340 1095.190 2028.400 ;
        RECT 1094.425 2028.200 1095.190 2028.340 ;
        RECT 1094.425 2028.155 1094.715 2028.200 ;
        RECT 1094.870 2028.140 1095.190 2028.200 ;
        RECT 1094.410 1980.400 1094.730 1980.460 ;
        RECT 1094.215 1980.260 1094.730 1980.400 ;
        RECT 1094.410 1980.200 1094.730 1980.260 ;
        RECT 1094.870 1863.100 1095.190 1863.160 ;
        RECT 1095.790 1863.100 1096.110 1863.160 ;
        RECT 1094.870 1862.960 1096.110 1863.100 ;
        RECT 1094.870 1862.900 1095.190 1862.960 ;
        RECT 1095.790 1862.900 1096.110 1862.960 ;
        RECT 1094.870 1838.960 1095.190 1839.020 ;
        RECT 1095.790 1838.960 1096.110 1839.020 ;
        RECT 1094.870 1838.820 1096.110 1838.960 ;
        RECT 1094.870 1838.760 1095.190 1838.820 ;
        RECT 1095.790 1838.760 1096.110 1838.820 ;
        RECT 1093.965 1801.220 1094.255 1801.265 ;
        RECT 1094.870 1801.220 1095.190 1801.280 ;
        RECT 1093.965 1801.080 1095.190 1801.220 ;
        RECT 1093.965 1801.035 1094.255 1801.080 ;
        RECT 1094.870 1801.020 1095.190 1801.080 ;
        RECT 1093.950 1774.020 1094.270 1774.080 ;
        RECT 1093.755 1773.880 1094.270 1774.020 ;
        RECT 1093.950 1773.820 1094.270 1773.880 ;
        RECT 1093.950 1773.340 1094.270 1773.400 ;
        RECT 1094.885 1773.340 1095.175 1773.385 ;
        RECT 1093.950 1773.200 1095.175 1773.340 ;
        RECT 1093.950 1773.140 1094.270 1773.200 ;
        RECT 1094.885 1773.155 1095.175 1773.200 ;
        RECT 1094.870 1752.260 1095.190 1752.320 ;
        RECT 1094.675 1752.120 1095.190 1752.260 ;
        RECT 1094.870 1752.060 1095.190 1752.120 ;
        RECT 1094.870 1704.660 1095.190 1704.720 ;
        RECT 1094.500 1704.520 1095.190 1704.660 ;
        RECT 1094.500 1704.380 1094.640 1704.520 ;
        RECT 1094.870 1704.460 1095.190 1704.520 ;
        RECT 1094.410 1704.120 1094.730 1704.380 ;
        RECT 1094.410 1689.020 1094.730 1689.080 ;
        RECT 1516.230 1689.020 1516.550 1689.080 ;
        RECT 1094.410 1688.880 1516.550 1689.020 ;
        RECT 1094.410 1688.820 1094.730 1688.880 ;
        RECT 1516.230 1688.820 1516.550 1688.880 ;
      LAYER via ;
        RECT 1094.900 3470.760 1095.160 3471.020 ;
        RECT 1095.820 3470.760 1096.080 3471.020 ;
        RECT 1095.820 3443.220 1096.080 3443.480 ;
        RECT 1095.360 3442.880 1095.620 3443.140 ;
        RECT 1094.900 3380.660 1095.160 3380.920 ;
        RECT 1095.360 3332.720 1095.620 3332.980 ;
        RECT 1095.820 3298.040 1096.080 3298.300 ;
        RECT 1096.740 3298.040 1097.000 3298.300 ;
        RECT 1096.740 3284.100 1097.000 3284.360 ;
        RECT 1096.280 3236.160 1096.540 3236.420 ;
        RECT 1096.280 3201.820 1096.540 3202.080 ;
        RECT 1095.360 3201.140 1095.620 3201.400 ;
        RECT 1095.360 3187.540 1095.620 3187.800 ;
        RECT 1095.820 3187.540 1096.080 3187.800 ;
        RECT 1096.740 3132.460 1097.000 3132.720 ;
        RECT 1096.740 3084.180 1097.000 3084.440 ;
        RECT 1096.740 3056.980 1097.000 3057.240 ;
        RECT 1095.360 3043.380 1095.620 3043.640 ;
        RECT 1095.360 3042.700 1095.620 3042.960 ;
        RECT 1096.280 3007.680 1096.540 3007.940 ;
        RECT 1096.280 2994.420 1096.540 2994.680 ;
        RECT 1095.820 2946.480 1096.080 2946.740 ;
        RECT 1094.900 2911.800 1095.160 2912.060 ;
        RECT 1095.820 2911.800 1096.080 2912.060 ;
        RECT 1094.900 2897.860 1095.160 2898.120 ;
        RECT 1094.440 2849.580 1094.700 2849.840 ;
        RECT 1094.440 2815.240 1094.700 2815.500 ;
        RECT 1094.900 2814.560 1095.160 2814.820 ;
        RECT 1094.440 2766.960 1094.700 2767.220 ;
        RECT 1094.440 2753.020 1094.700 2753.280 ;
        RECT 1094.440 2718.680 1094.700 2718.940 ;
        RECT 1094.900 2718.000 1095.160 2718.260 ;
        RECT 1094.900 2621.440 1095.160 2621.700 ;
        RECT 1095.820 2621.440 1096.080 2621.700 ;
        RECT 1094.440 2511.620 1094.700 2511.880 ;
        RECT 1096.740 2511.620 1097.000 2511.880 ;
        RECT 1095.820 2401.120 1096.080 2401.380 ;
        RECT 1096.740 2401.120 1097.000 2401.380 ;
        RECT 1095.820 2304.560 1096.080 2304.820 ;
        RECT 1096.740 2304.560 1097.000 2304.820 ;
        RECT 1096.280 2221.600 1096.540 2221.860 ;
        RECT 1097.200 2221.600 1097.460 2221.860 ;
        RECT 1094.900 2138.980 1095.160 2139.240 ;
        RECT 1095.820 2138.980 1096.080 2139.240 ;
        RECT 1093.520 2125.040 1093.780 2125.300 ;
        RECT 1094.900 2125.040 1095.160 2125.300 ;
        RECT 1094.440 2042.420 1094.700 2042.680 ;
        RECT 1094.900 2041.740 1095.160 2042.000 ;
        RECT 1094.900 2028.140 1095.160 2028.400 ;
        RECT 1094.440 1980.200 1094.700 1980.460 ;
        RECT 1094.900 1862.900 1095.160 1863.160 ;
        RECT 1095.820 1862.900 1096.080 1863.160 ;
        RECT 1094.900 1838.760 1095.160 1839.020 ;
        RECT 1095.820 1838.760 1096.080 1839.020 ;
        RECT 1094.900 1801.020 1095.160 1801.280 ;
        RECT 1093.980 1773.820 1094.240 1774.080 ;
        RECT 1093.980 1773.140 1094.240 1773.400 ;
        RECT 1094.900 1752.060 1095.160 1752.320 ;
        RECT 1094.900 1704.460 1095.160 1704.720 ;
        RECT 1094.440 1704.120 1094.700 1704.380 ;
        RECT 1094.440 1688.820 1094.700 1689.080 ;
        RECT 1516.260 1688.820 1516.520 1689.080 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3471.050 1095.100 3517.600 ;
        RECT 1094.900 3470.730 1095.160 3471.050 ;
        RECT 1095.820 3470.730 1096.080 3471.050 ;
        RECT 1095.880 3443.510 1096.020 3470.730 ;
        RECT 1095.820 3443.190 1096.080 3443.510 ;
        RECT 1095.360 3442.850 1095.620 3443.170 ;
        RECT 1095.420 3394.970 1095.560 3442.850 ;
        RECT 1094.960 3394.830 1095.560 3394.970 ;
        RECT 1094.960 3380.950 1095.100 3394.830 ;
        RECT 1094.900 3380.630 1095.160 3380.950 ;
        RECT 1095.360 3332.690 1095.620 3333.010 ;
        RECT 1095.420 3298.410 1095.560 3332.690 ;
        RECT 1095.420 3298.330 1096.020 3298.410 ;
        RECT 1095.420 3298.270 1096.080 3298.330 ;
        RECT 1095.820 3298.010 1096.080 3298.270 ;
        RECT 1096.740 3298.010 1097.000 3298.330 ;
        RECT 1096.800 3284.390 1096.940 3298.010 ;
        RECT 1096.740 3284.070 1097.000 3284.390 ;
        RECT 1096.280 3236.130 1096.540 3236.450 ;
        RECT 1096.340 3202.110 1096.480 3236.130 ;
        RECT 1096.280 3201.790 1096.540 3202.110 ;
        RECT 1095.360 3201.110 1095.620 3201.430 ;
        RECT 1095.420 3187.830 1095.560 3201.110 ;
        RECT 1095.360 3187.510 1095.620 3187.830 ;
        RECT 1095.820 3187.510 1096.080 3187.830 ;
        RECT 1095.880 3152.890 1096.020 3187.510 ;
        RECT 1095.880 3152.750 1096.940 3152.890 ;
        RECT 1096.800 3132.750 1096.940 3152.750 ;
        RECT 1096.740 3132.430 1097.000 3132.750 ;
        RECT 1096.740 3084.150 1097.000 3084.470 ;
        RECT 1096.800 3057.270 1096.940 3084.150 ;
        RECT 1096.740 3056.950 1097.000 3057.270 ;
        RECT 1095.360 3043.350 1095.620 3043.670 ;
        RECT 1095.420 3042.990 1095.560 3043.350 ;
        RECT 1095.360 3042.670 1095.620 3042.990 ;
        RECT 1096.280 3007.650 1096.540 3007.970 ;
        RECT 1096.340 2994.710 1096.480 3007.650 ;
        RECT 1096.280 2994.390 1096.540 2994.710 ;
        RECT 1095.820 2946.450 1096.080 2946.770 ;
        RECT 1095.880 2912.090 1096.020 2946.450 ;
        RECT 1094.900 2911.770 1095.160 2912.090 ;
        RECT 1095.820 2911.770 1096.080 2912.090 ;
        RECT 1094.960 2898.150 1095.100 2911.770 ;
        RECT 1094.900 2897.830 1095.160 2898.150 ;
        RECT 1094.440 2849.550 1094.700 2849.870 ;
        RECT 1094.500 2815.530 1094.640 2849.550 ;
        RECT 1094.440 2815.210 1094.700 2815.530 ;
        RECT 1094.900 2814.530 1095.160 2814.850 ;
        RECT 1094.960 2801.330 1095.100 2814.530 ;
        RECT 1094.500 2801.190 1095.100 2801.330 ;
        RECT 1094.500 2767.250 1094.640 2801.190 ;
        RECT 1094.440 2766.930 1094.700 2767.250 ;
        RECT 1094.440 2752.990 1094.700 2753.310 ;
        RECT 1094.500 2718.970 1094.640 2752.990 ;
        RECT 1094.440 2718.650 1094.700 2718.970 ;
        RECT 1094.900 2717.970 1095.160 2718.290 ;
        RECT 1094.960 2704.885 1095.100 2717.970 ;
        RECT 1094.890 2704.515 1095.170 2704.885 ;
        RECT 1095.810 2704.515 1096.090 2704.885 ;
        RECT 1095.880 2669.410 1096.020 2704.515 ;
        RECT 1094.960 2669.270 1096.020 2669.410 ;
        RECT 1094.960 2656.605 1095.100 2669.270 ;
        RECT 1094.890 2656.235 1095.170 2656.605 ;
        RECT 1095.810 2656.235 1096.090 2656.605 ;
        RECT 1095.880 2621.730 1096.020 2656.235 ;
        RECT 1094.900 2621.410 1095.160 2621.730 ;
        RECT 1095.820 2621.410 1096.080 2621.730 ;
        RECT 1094.960 2573.530 1095.100 2621.410 ;
        RECT 1094.960 2573.390 1095.560 2573.530 ;
        RECT 1095.420 2560.045 1095.560 2573.390 ;
        RECT 1094.430 2559.675 1094.710 2560.045 ;
        RECT 1095.350 2559.675 1095.630 2560.045 ;
        RECT 1094.500 2511.910 1094.640 2559.675 ;
        RECT 1094.440 2511.590 1094.700 2511.910 ;
        RECT 1096.740 2511.590 1097.000 2511.910 ;
        RECT 1096.800 2476.970 1096.940 2511.590 ;
        RECT 1096.340 2476.830 1096.940 2476.970 ;
        RECT 1096.340 2429.370 1096.480 2476.830 ;
        RECT 1095.880 2429.230 1096.480 2429.370 ;
        RECT 1095.880 2401.410 1096.020 2429.230 ;
        RECT 1095.820 2401.090 1096.080 2401.410 ;
        RECT 1096.740 2401.090 1097.000 2401.410 ;
        RECT 1096.800 2400.810 1096.940 2401.090 ;
        RECT 1096.340 2400.670 1096.940 2400.810 ;
        RECT 1096.340 2353.210 1096.480 2400.670 ;
        RECT 1095.880 2353.070 1096.480 2353.210 ;
        RECT 1095.880 2304.850 1096.020 2353.070 ;
        RECT 1095.820 2304.530 1096.080 2304.850 ;
        RECT 1096.740 2304.530 1097.000 2304.850 ;
        RECT 1096.800 2304.250 1096.940 2304.530 ;
        RECT 1096.340 2304.110 1096.940 2304.250 ;
        RECT 1096.340 2221.890 1096.480 2304.110 ;
        RECT 1096.280 2221.570 1096.540 2221.890 ;
        RECT 1097.200 2221.570 1097.460 2221.890 ;
        RECT 1097.260 2173.805 1097.400 2221.570 ;
        RECT 1095.810 2173.435 1096.090 2173.805 ;
        RECT 1097.190 2173.435 1097.470 2173.805 ;
        RECT 1095.880 2139.270 1096.020 2173.435 ;
        RECT 1094.900 2138.950 1095.160 2139.270 ;
        RECT 1095.820 2138.950 1096.080 2139.270 ;
        RECT 1094.960 2125.330 1095.100 2138.950 ;
        RECT 1093.520 2125.010 1093.780 2125.330 ;
        RECT 1094.900 2125.010 1095.160 2125.330 ;
        RECT 1093.580 2077.245 1093.720 2125.010 ;
        RECT 1093.510 2076.875 1093.790 2077.245 ;
        RECT 1094.430 2076.875 1094.710 2077.245 ;
        RECT 1094.500 2042.710 1094.640 2076.875 ;
        RECT 1094.440 2042.390 1094.700 2042.710 ;
        RECT 1094.900 2041.710 1095.160 2042.030 ;
        RECT 1094.960 2028.430 1095.100 2041.710 ;
        RECT 1094.900 2028.110 1095.160 2028.430 ;
        RECT 1094.440 1980.170 1094.700 1980.490 ;
        RECT 1094.500 1979.890 1094.640 1980.170 ;
        RECT 1094.040 1979.750 1094.640 1979.890 ;
        RECT 1094.040 1945.210 1094.180 1979.750 ;
        RECT 1094.040 1945.070 1095.100 1945.210 ;
        RECT 1094.960 1863.190 1095.100 1945.070 ;
        RECT 1094.900 1862.870 1095.160 1863.190 ;
        RECT 1095.820 1862.870 1096.080 1863.190 ;
        RECT 1095.880 1839.050 1096.020 1862.870 ;
        RECT 1094.900 1838.730 1095.160 1839.050 ;
        RECT 1095.820 1838.730 1096.080 1839.050 ;
        RECT 1094.960 1801.310 1095.100 1838.730 ;
        RECT 1094.900 1800.990 1095.160 1801.310 ;
        RECT 1093.980 1773.790 1094.240 1774.110 ;
        RECT 1094.040 1773.430 1094.180 1773.790 ;
        RECT 1093.980 1773.110 1094.240 1773.430 ;
        RECT 1094.900 1752.030 1095.160 1752.350 ;
        RECT 1094.960 1704.750 1095.100 1752.030 ;
        RECT 1094.900 1704.430 1095.160 1704.750 ;
        RECT 1094.440 1704.090 1094.700 1704.410 ;
        RECT 1094.500 1689.110 1094.640 1704.090 ;
        RECT 1516.330 1700.340 1516.610 1704.000 ;
        RECT 1516.320 1700.000 1516.610 1700.340 ;
        RECT 1516.320 1689.110 1516.460 1700.000 ;
        RECT 1094.440 1688.790 1094.700 1689.110 ;
        RECT 1516.260 1688.790 1516.520 1689.110 ;
      LAYER via2 ;
        RECT 1094.890 2704.560 1095.170 2704.840 ;
        RECT 1095.810 2704.560 1096.090 2704.840 ;
        RECT 1094.890 2656.280 1095.170 2656.560 ;
        RECT 1095.810 2656.280 1096.090 2656.560 ;
        RECT 1094.430 2559.720 1094.710 2560.000 ;
        RECT 1095.350 2559.720 1095.630 2560.000 ;
        RECT 1095.810 2173.480 1096.090 2173.760 ;
        RECT 1097.190 2173.480 1097.470 2173.760 ;
        RECT 1093.510 2076.920 1093.790 2077.200 ;
        RECT 1094.430 2076.920 1094.710 2077.200 ;
      LAYER met3 ;
        RECT 1094.865 2704.850 1095.195 2704.865 ;
        RECT 1095.785 2704.850 1096.115 2704.865 ;
        RECT 1094.865 2704.550 1096.115 2704.850 ;
        RECT 1094.865 2704.535 1095.195 2704.550 ;
        RECT 1095.785 2704.535 1096.115 2704.550 ;
        RECT 1094.865 2656.570 1095.195 2656.585 ;
        RECT 1095.785 2656.570 1096.115 2656.585 ;
        RECT 1094.865 2656.270 1096.115 2656.570 ;
        RECT 1094.865 2656.255 1095.195 2656.270 ;
        RECT 1095.785 2656.255 1096.115 2656.270 ;
        RECT 1094.405 2560.010 1094.735 2560.025 ;
        RECT 1095.325 2560.010 1095.655 2560.025 ;
        RECT 1094.405 2559.710 1095.655 2560.010 ;
        RECT 1094.405 2559.695 1094.735 2559.710 ;
        RECT 1095.325 2559.695 1095.655 2559.710 ;
        RECT 1095.785 2173.770 1096.115 2173.785 ;
        RECT 1097.165 2173.770 1097.495 2173.785 ;
        RECT 1095.785 2173.470 1097.495 2173.770 ;
        RECT 1095.785 2173.455 1096.115 2173.470 ;
        RECT 1097.165 2173.455 1097.495 2173.470 ;
        RECT 1093.485 2077.210 1093.815 2077.225 ;
        RECT 1094.405 2077.210 1094.735 2077.225 ;
        RECT 1093.485 2076.910 1094.735 2077.210 ;
        RECT 1093.485 2076.895 1093.815 2076.910 ;
        RECT 1094.405 2076.895 1094.735 2076.910 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
        RECT 771.565 2898.585 771.735 2946.355 ;
        RECT 772.025 2608.225 772.195 2656.335 ;
        RECT 772.025 2511.665 772.195 2559.775 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
        RECT 771.565 2946.185 771.735 2946.355 ;
        RECT 772.025 2656.165 772.195 2656.335 ;
        RECT 772.025 2559.605 772.195 2559.775 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 771.490 3174.140 771.810 3174.200 ;
        RECT 772.410 3174.140 772.730 3174.200 ;
        RECT 771.490 3174.000 772.730 3174.140 ;
        RECT 771.490 3173.940 771.810 3174.000 ;
        RECT 772.410 3173.940 772.730 3174.000 ;
        RECT 771.490 3077.580 771.810 3077.640 ;
        RECT 772.410 3077.580 772.730 3077.640 ;
        RECT 771.490 3077.440 772.730 3077.580 ;
        RECT 771.490 3077.380 771.810 3077.440 ;
        RECT 772.410 3077.380 772.730 3077.440 ;
        RECT 771.490 2981.020 771.810 2981.080 ;
        RECT 772.410 2981.020 772.730 2981.080 ;
        RECT 771.490 2980.880 772.730 2981.020 ;
        RECT 771.490 2980.820 771.810 2980.880 ;
        RECT 772.410 2980.820 772.730 2980.880 ;
        RECT 771.490 2946.340 771.810 2946.400 ;
        RECT 771.295 2946.200 771.810 2946.340 ;
        RECT 771.490 2946.140 771.810 2946.200 ;
        RECT 771.490 2898.740 771.810 2898.800 ;
        RECT 771.295 2898.600 771.810 2898.740 ;
        RECT 771.490 2898.540 771.810 2898.600 ;
        RECT 771.030 2898.060 771.350 2898.120 ;
        RECT 771.950 2898.060 772.270 2898.120 ;
        RECT 771.030 2897.920 772.270 2898.060 ;
        RECT 771.030 2897.860 771.350 2897.920 ;
        RECT 771.950 2897.860 772.270 2897.920 ;
        RECT 771.030 2814.760 771.350 2814.820 ;
        RECT 771.950 2814.760 772.270 2814.820 ;
        RECT 771.030 2814.620 772.270 2814.760 ;
        RECT 771.030 2814.560 771.350 2814.620 ;
        RECT 771.950 2814.560 772.270 2814.620 ;
        RECT 771.950 2656.320 772.270 2656.380 ;
        RECT 771.755 2656.180 772.270 2656.320 ;
        RECT 771.950 2656.120 772.270 2656.180 ;
        RECT 771.965 2608.380 772.255 2608.425 ;
        RECT 772.410 2608.380 772.730 2608.440 ;
        RECT 771.965 2608.240 772.730 2608.380 ;
        RECT 771.965 2608.195 772.255 2608.240 ;
        RECT 772.410 2608.180 772.730 2608.240 ;
        RECT 771.950 2559.760 772.270 2559.820 ;
        RECT 771.755 2559.620 772.270 2559.760 ;
        RECT 771.950 2559.560 772.270 2559.620 ;
        RECT 771.965 2511.820 772.255 2511.865 ;
        RECT 772.410 2511.820 772.730 2511.880 ;
        RECT 771.965 2511.680 772.730 2511.820 ;
        RECT 771.965 2511.635 772.255 2511.680 ;
        RECT 772.410 2511.620 772.730 2511.680 ;
        RECT 771.490 2429.000 771.810 2429.260 ;
        RECT 771.580 2428.520 771.720 2429.000 ;
        RECT 771.950 2428.520 772.270 2428.580 ;
        RECT 771.580 2428.380 772.270 2428.520 ;
        RECT 771.950 2428.320 772.270 2428.380 ;
        RECT 770.570 2414.920 770.890 2414.980 ;
        RECT 771.950 2414.920 772.270 2414.980 ;
        RECT 770.570 2414.780 772.270 2414.920 ;
        RECT 770.570 2414.720 770.890 2414.780 ;
        RECT 771.950 2414.720 772.270 2414.780 ;
        RECT 771.490 2363.240 771.810 2363.300 ;
        RECT 1382.370 2363.240 1382.690 2363.300 ;
        RECT 771.490 2363.100 1382.690 2363.240 ;
        RECT 771.490 2363.040 771.810 2363.100 ;
        RECT 1382.370 2363.040 1382.690 2363.100 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 771.520 3173.940 771.780 3174.200 ;
        RECT 772.440 3173.940 772.700 3174.200 ;
        RECT 771.520 3077.380 771.780 3077.640 ;
        RECT 772.440 3077.380 772.700 3077.640 ;
        RECT 771.520 2980.820 771.780 2981.080 ;
        RECT 772.440 2980.820 772.700 2981.080 ;
        RECT 771.520 2946.140 771.780 2946.400 ;
        RECT 771.520 2898.540 771.780 2898.800 ;
        RECT 771.060 2897.860 771.320 2898.120 ;
        RECT 771.980 2897.860 772.240 2898.120 ;
        RECT 771.060 2814.560 771.320 2814.820 ;
        RECT 771.980 2814.560 772.240 2814.820 ;
        RECT 771.980 2656.120 772.240 2656.380 ;
        RECT 772.440 2608.180 772.700 2608.440 ;
        RECT 771.980 2559.560 772.240 2559.820 ;
        RECT 772.440 2511.620 772.700 2511.880 ;
        RECT 771.520 2429.000 771.780 2429.260 ;
        RECT 771.980 2428.320 772.240 2428.580 ;
        RECT 770.600 2414.720 770.860 2414.980 ;
        RECT 771.980 2414.720 772.240 2414.980 ;
        RECT 771.520 2363.040 771.780 2363.300 ;
        RECT 1382.400 2363.040 1382.660 2363.300 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3222.250 772.640 3270.470 ;
        RECT 771.580 3222.110 772.640 3222.250 ;
        RECT 771.580 3174.230 771.720 3222.110 ;
        RECT 771.520 3173.910 771.780 3174.230 ;
        RECT 772.440 3173.910 772.700 3174.230 ;
        RECT 772.500 3125.690 772.640 3173.910 ;
        RECT 771.580 3125.550 772.640 3125.690 ;
        RECT 771.580 3077.670 771.720 3125.550 ;
        RECT 771.520 3077.350 771.780 3077.670 ;
        RECT 772.440 3077.350 772.700 3077.670 ;
        RECT 772.500 3029.130 772.640 3077.350 ;
        RECT 771.580 3028.990 772.640 3029.130 ;
        RECT 771.580 2981.110 771.720 3028.990 ;
        RECT 771.520 2980.790 771.780 2981.110 ;
        RECT 772.440 2980.850 772.700 2981.110 ;
        RECT 772.040 2980.790 772.700 2980.850 ;
        RECT 772.040 2980.710 772.640 2980.790 ;
        RECT 772.040 2959.770 772.180 2980.710 ;
        RECT 771.580 2959.630 772.180 2959.770 ;
        RECT 771.580 2946.430 771.720 2959.630 ;
        RECT 771.520 2946.110 771.780 2946.430 ;
        RECT 771.520 2898.570 771.780 2898.830 ;
        RECT 771.120 2898.510 771.780 2898.570 ;
        RECT 771.120 2898.430 771.720 2898.510 ;
        RECT 771.120 2898.150 771.260 2898.430 ;
        RECT 771.060 2897.830 771.320 2898.150 ;
        RECT 771.980 2897.830 772.240 2898.150 ;
        RECT 772.040 2814.850 772.180 2897.830 ;
        RECT 771.060 2814.530 771.320 2814.850 ;
        RECT 771.980 2814.530 772.240 2814.850 ;
        RECT 771.120 2766.650 771.260 2814.530 ;
        RECT 771.120 2766.510 771.720 2766.650 ;
        RECT 771.580 2719.050 771.720 2766.510 ;
        RECT 771.580 2718.910 772.640 2719.050 ;
        RECT 772.500 2670.090 772.640 2718.910 ;
        RECT 772.040 2669.950 772.640 2670.090 ;
        RECT 772.040 2656.410 772.180 2669.950 ;
        RECT 771.980 2656.090 772.240 2656.410 ;
        RECT 772.440 2608.150 772.700 2608.470 ;
        RECT 772.500 2573.530 772.640 2608.150 ;
        RECT 772.040 2573.390 772.640 2573.530 ;
        RECT 772.040 2559.850 772.180 2573.390 ;
        RECT 771.980 2559.530 772.240 2559.850 ;
        RECT 772.440 2511.590 772.700 2511.910 ;
        RECT 772.500 2476.970 772.640 2511.590 ;
        RECT 771.580 2476.830 772.640 2476.970 ;
        RECT 771.580 2429.290 771.720 2476.830 ;
        RECT 771.520 2428.970 771.780 2429.290 ;
        RECT 771.980 2428.290 772.240 2428.610 ;
        RECT 772.040 2415.010 772.180 2428.290 ;
        RECT 770.600 2414.690 770.860 2415.010 ;
        RECT 771.980 2414.690 772.240 2415.010 ;
        RECT 770.660 2366.925 770.800 2414.690 ;
        RECT 770.590 2366.555 770.870 2366.925 ;
        RECT 771.510 2366.555 771.790 2366.925 ;
        RECT 771.580 2363.330 771.720 2366.555 ;
        RECT 771.520 2363.010 771.780 2363.330 ;
        RECT 1382.400 2363.010 1382.660 2363.330 ;
        RECT 1382.460 2350.000 1382.600 2363.010 ;
        RECT 1382.460 2349.740 1382.750 2350.000 ;
        RECT 1382.470 2346.000 1382.750 2349.740 ;
      LAYER via2 ;
        RECT 770.590 2366.600 770.870 2366.880 ;
        RECT 771.510 2366.600 771.790 2366.880 ;
      LAYER met3 ;
        RECT 770.565 2366.890 770.895 2366.905 ;
        RECT 771.485 2366.890 771.815 2366.905 ;
        RECT 770.565 2366.590 771.815 2366.890 ;
        RECT 770.565 2366.575 770.895 2366.590 ;
        RECT 771.485 2366.575 771.815 2366.590 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1794.070 3501.560 1794.390 3501.620 ;
        RECT 121.510 3501.420 1794.390 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1794.070 3501.360 1794.390 3501.420 ;
        RECT 1795.910 2028.000 1796.230 2028.060 ;
        RECT 1797.750 2028.000 1798.070 2028.060 ;
        RECT 1795.910 2027.860 1798.070 2028.000 ;
        RECT 1795.910 2027.800 1796.230 2027.860 ;
        RECT 1797.750 2027.800 1798.070 2027.860 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1794.100 3501.360 1794.360 3501.620 ;
        RECT 1795.940 2027.800 1796.200 2028.060 ;
        RECT 1797.780 2027.800 1798.040 2028.060 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1794.100 3501.330 1794.360 3501.650 ;
        RECT 1794.160 2028.170 1794.300 3501.330 ;
        RECT 1794.160 2028.090 1796.140 2028.170 ;
        RECT 1794.160 2028.030 1796.200 2028.090 ;
        RECT 1795.940 2027.770 1796.200 2028.030 ;
        RECT 1797.780 2027.770 1798.040 2028.090 ;
        RECT 1797.840 2027.605 1797.980 2027.770 ;
        RECT 1797.770 2027.235 1798.050 2027.605 ;
      LAYER via2 ;
        RECT 1797.770 2027.280 1798.050 2027.560 ;
      LAYER met3 ;
        RECT 1797.745 2027.570 1798.075 2027.585 ;
        RECT 1797.745 2027.255 1798.290 2027.570 ;
        RECT 1797.990 2025.000 1798.290 2027.255 ;
        RECT 1797.000 2024.400 1801.000 2025.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1690.040 17.410 1690.100 ;
        RECT 1353.850 1690.040 1354.170 1690.100 ;
        RECT 17.090 1689.900 1354.170 1690.040 ;
        RECT 17.090 1689.840 17.410 1689.900 ;
        RECT 1353.850 1689.840 1354.170 1689.900 ;
      LAYER via ;
        RECT 17.120 1689.840 17.380 1690.100 ;
        RECT 1353.880 1689.840 1354.140 1690.100 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 1690.130 17.320 3339.635 ;
        RECT 1353.950 1700.340 1354.230 1704.000 ;
        RECT 1353.940 1700.000 1354.230 1700.340 ;
        RECT 1353.940 1690.130 1354.080 1700.000 ;
        RECT 17.120 1689.810 17.380 1690.130 ;
        RECT 1353.880 1689.810 1354.140 1690.130 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2477.480 16.950 2477.540 ;
        RECT 1795.450 2477.480 1795.770 2477.540 ;
        RECT 16.630 2477.340 1795.770 2477.480 ;
        RECT 16.630 2477.280 16.950 2477.340 ;
        RECT 1795.450 2477.280 1795.770 2477.340 ;
      LAYER via ;
        RECT 16.660 2477.280 16.920 2477.540 ;
        RECT 1795.480 2477.280 1795.740 2477.540 ;
      LAYER met2 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 16.660 2477.250 16.920 2477.395 ;
        RECT 1795.480 2477.250 1795.740 2477.570 ;
        RECT 1795.540 2315.810 1795.680 2477.250 ;
        RECT 1797.770 2315.810 1798.050 2315.925 ;
        RECT 1795.540 2315.670 1798.050 2315.810 ;
        RECT 1797.770 2315.555 1798.050 2315.670 ;
      LAYER via2 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
        RECT 1797.770 2315.600 1798.050 2315.880 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
        RECT 1797.745 2315.890 1798.075 2315.905 ;
        RECT 1797.745 2315.575 1798.290 2315.890 ;
        RECT 1797.990 2314.000 1798.290 2315.575 ;
        RECT 1797.000 2313.400 1801.000 2314.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2360.180 18.790 2360.240 ;
        RECT 1754.050 2360.180 1754.370 2360.240 ;
        RECT 18.470 2360.040 1754.370 2360.180 ;
        RECT 18.470 2359.980 18.790 2360.040 ;
        RECT 1754.050 2359.980 1754.370 2360.040 ;
      LAYER via ;
        RECT 18.500 2359.980 18.760 2360.240 ;
        RECT 1754.080 2359.980 1754.340 2360.240 ;
      LAYER met2 ;
        RECT 18.500 2359.950 18.760 2360.270 ;
        RECT 1754.080 2359.950 1754.340 2360.270 ;
        RECT 18.560 2190.125 18.700 2359.950 ;
        RECT 1754.140 2350.000 1754.280 2359.950 ;
        RECT 1754.140 2349.740 1754.430 2350.000 ;
        RECT 1754.150 2346.000 1754.430 2349.740 ;
        RECT 18.490 2189.755 18.770 2190.125 ;
      LAYER via2 ;
        RECT 18.490 2189.800 18.770 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 18.465 2190.090 18.795 2190.105 ;
        RECT -4.800 2189.790 18.795 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 18.465 2189.775 18.795 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 1686.980 18.790 1687.040 ;
        RECT 1678.610 1686.980 1678.930 1687.040 ;
        RECT 18.470 1686.840 1678.930 1686.980 ;
        RECT 18.470 1686.780 18.790 1686.840 ;
        RECT 1678.610 1686.780 1678.930 1686.840 ;
      LAYER via ;
        RECT 18.500 1686.780 18.760 1687.040 ;
        RECT 1678.640 1686.780 1678.900 1687.040 ;
      LAYER met2 ;
        RECT 1678.710 1700.340 1678.990 1704.000 ;
        RECT 1678.700 1700.000 1678.990 1700.340 ;
        RECT 1678.700 1687.070 1678.840 1700.000 ;
        RECT 18.500 1686.750 18.760 1687.070 ;
        RECT 1678.640 1686.750 1678.900 1687.070 ;
        RECT 18.560 1615.525 18.700 1686.750 ;
        RECT 18.490 1615.155 18.770 1615.525 ;
      LAYER via2 ;
        RECT 18.490 1615.200 18.770 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 18.465 1615.490 18.795 1615.505 ;
        RECT -4.800 1615.190 18.795 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 18.465 1615.175 18.795 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1795.910 1947.420 1796.230 1947.480 ;
        RECT 1797.750 1947.420 1798.070 1947.480 ;
        RECT 1795.910 1947.280 1798.070 1947.420 ;
        RECT 1795.910 1947.220 1796.230 1947.280 ;
        RECT 1797.750 1947.220 1798.070 1947.280 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 1794.530 1400.700 1794.850 1400.760 ;
        RECT 17.090 1400.560 1794.850 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 1794.530 1400.500 1794.850 1400.560 ;
      LAYER via ;
        RECT 1795.940 1947.220 1796.200 1947.480 ;
        RECT 1797.780 1947.220 1798.040 1947.480 ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 1794.560 1400.500 1794.820 1400.760 ;
      LAYER met2 ;
        RECT 1797.770 1949.715 1798.050 1950.085 ;
        RECT 1797.840 1947.510 1797.980 1949.715 ;
        RECT 1795.940 1947.250 1796.200 1947.510 ;
        RECT 1795.080 1947.190 1796.200 1947.250 ;
        RECT 1797.780 1947.190 1798.040 1947.510 ;
        RECT 1795.080 1947.110 1796.140 1947.190 ;
        RECT 1795.080 1942.490 1795.220 1947.110 ;
        RECT 1794.620 1942.350 1795.220 1942.490 ;
        RECT 1794.620 1896.930 1794.760 1942.350 ;
        RECT 1794.620 1896.790 1795.220 1896.930 ;
        RECT 1795.080 1849.330 1795.220 1896.790 ;
        RECT 1795.080 1849.190 1795.680 1849.330 ;
        RECT 1795.540 1821.960 1795.680 1849.190 ;
        RECT 1794.620 1821.820 1795.680 1821.960 ;
        RECT 1794.620 1773.170 1794.760 1821.820 ;
        RECT 1794.160 1773.030 1794.760 1773.170 ;
        RECT 1794.160 1758.890 1794.300 1773.030 ;
        RECT 1793.700 1758.750 1794.300 1758.890 ;
        RECT 1793.700 1752.090 1793.840 1758.750 ;
        RECT 1793.700 1751.950 1794.760 1752.090 ;
        RECT 1794.620 1400.790 1794.760 1751.950 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 1794.560 1400.470 1794.820 1400.790 ;
      LAYER via2 ;
        RECT 1797.770 1949.760 1798.050 1950.040 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 1797.000 1952.320 1801.000 1952.920 ;
        RECT 1797.990 1950.065 1798.290 1952.320 ;
        RECT 1797.745 1949.750 1798.290 1950.065 ;
        RECT 1797.745 1949.735 1798.075 1949.750 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1796.445 1800.385 1796.615 1828.435 ;
        RECT 1794.145 1256.045 1794.315 1304.155 ;
        RECT 1794.605 1173.085 1794.775 1207.255 ;
      LAYER mcon ;
        RECT 1796.445 1828.265 1796.615 1828.435 ;
        RECT 1794.145 1303.985 1794.315 1304.155 ;
        RECT 1794.605 1207.085 1794.775 1207.255 ;
      LAYER met1 ;
        RECT 1796.370 1877.040 1796.690 1877.100 ;
        RECT 1797.750 1877.040 1798.070 1877.100 ;
        RECT 1796.370 1876.900 1798.070 1877.040 ;
        RECT 1796.370 1876.840 1796.690 1876.900 ;
        RECT 1797.750 1876.840 1798.070 1876.900 ;
        RECT 1796.370 1828.420 1796.690 1828.480 ;
        RECT 1796.175 1828.280 1796.690 1828.420 ;
        RECT 1796.370 1828.220 1796.690 1828.280 ;
        RECT 1795.910 1800.540 1796.230 1800.600 ;
        RECT 1796.385 1800.540 1796.675 1800.585 ;
        RECT 1795.910 1800.400 1796.675 1800.540 ;
        RECT 1795.910 1800.340 1796.230 1800.400 ;
        RECT 1796.385 1800.355 1796.675 1800.400 ;
        RECT 1794.070 1676.780 1794.390 1676.840 ;
        RECT 1795.450 1676.780 1795.770 1676.840 ;
        RECT 1794.070 1676.640 1795.770 1676.780 ;
        RECT 1794.070 1676.580 1794.390 1676.640 ;
        RECT 1795.450 1676.580 1795.770 1676.640 ;
        RECT 1794.070 1628.160 1794.390 1628.220 ;
        RECT 1795.450 1628.160 1795.770 1628.220 ;
        RECT 1794.070 1628.020 1795.770 1628.160 ;
        RECT 1794.070 1627.960 1794.390 1628.020 ;
        RECT 1795.450 1627.960 1795.770 1628.020 ;
        RECT 1794.070 1580.220 1794.390 1580.280 ;
        RECT 1795.450 1580.220 1795.770 1580.280 ;
        RECT 1794.070 1580.080 1795.770 1580.220 ;
        RECT 1794.070 1580.020 1794.390 1580.080 ;
        RECT 1795.450 1580.020 1795.770 1580.080 ;
        RECT 1794.070 1531.600 1794.390 1531.660 ;
        RECT 1795.450 1531.600 1795.770 1531.660 ;
        RECT 1794.070 1531.460 1795.770 1531.600 ;
        RECT 1794.070 1531.400 1794.390 1531.460 ;
        RECT 1795.450 1531.400 1795.770 1531.460 ;
        RECT 1794.070 1483.660 1794.390 1483.720 ;
        RECT 1795.450 1483.660 1795.770 1483.720 ;
        RECT 1794.070 1483.520 1795.770 1483.660 ;
        RECT 1794.070 1483.460 1794.390 1483.520 ;
        RECT 1795.450 1483.460 1795.770 1483.520 ;
        RECT 1794.070 1435.040 1794.390 1435.100 ;
        RECT 1795.450 1435.040 1795.770 1435.100 ;
        RECT 1794.070 1434.900 1795.770 1435.040 ;
        RECT 1794.070 1434.840 1794.390 1434.900 ;
        RECT 1795.450 1434.840 1795.770 1434.900 ;
        RECT 1794.070 1387.100 1794.390 1387.160 ;
        RECT 1795.450 1387.100 1795.770 1387.160 ;
        RECT 1794.070 1386.960 1795.770 1387.100 ;
        RECT 1794.070 1386.900 1794.390 1386.960 ;
        RECT 1795.450 1386.900 1795.770 1386.960 ;
        RECT 1794.070 1338.820 1794.390 1338.880 ;
        RECT 1794.990 1338.820 1795.310 1338.880 ;
        RECT 1794.070 1338.680 1795.310 1338.820 ;
        RECT 1794.070 1338.620 1794.390 1338.680 ;
        RECT 1794.990 1338.620 1795.310 1338.680 ;
        RECT 1794.085 1304.140 1794.375 1304.185 ;
        RECT 1794.530 1304.140 1794.850 1304.200 ;
        RECT 1794.085 1304.000 1794.850 1304.140 ;
        RECT 1794.085 1303.955 1794.375 1304.000 ;
        RECT 1794.530 1303.940 1794.850 1304.000 ;
        RECT 1794.070 1256.200 1794.390 1256.260 ;
        RECT 1793.875 1256.060 1794.390 1256.200 ;
        RECT 1794.070 1256.000 1794.390 1256.060 ;
        RECT 1794.530 1207.240 1794.850 1207.300 ;
        RECT 1794.335 1207.100 1794.850 1207.240 ;
        RECT 1794.530 1207.040 1794.850 1207.100 ;
        RECT 1794.545 1173.240 1794.835 1173.285 ;
        RECT 1795.450 1173.240 1795.770 1173.300 ;
        RECT 1794.545 1173.100 1795.770 1173.240 ;
        RECT 1794.545 1173.055 1794.835 1173.100 ;
        RECT 1795.450 1173.040 1795.770 1173.100 ;
        RECT 1794.530 1111.020 1794.850 1111.080 ;
        RECT 1795.910 1111.020 1796.230 1111.080 ;
        RECT 1794.530 1110.880 1796.230 1111.020 ;
        RECT 1794.530 1110.820 1794.850 1110.880 ;
        RECT 1795.910 1110.820 1796.230 1110.880 ;
        RECT 1795.910 1077.020 1796.230 1077.080 ;
        RECT 1795.540 1076.880 1796.230 1077.020 ;
        RECT 1795.540 1076.400 1795.680 1076.880 ;
        RECT 1795.910 1076.820 1796.230 1076.880 ;
        RECT 1795.450 1076.140 1795.770 1076.400 ;
        RECT 1794.530 1014.460 1794.850 1014.520 ;
        RECT 1795.910 1014.460 1796.230 1014.520 ;
        RECT 1794.530 1014.320 1796.230 1014.460 ;
        RECT 1794.530 1014.260 1794.850 1014.320 ;
        RECT 1795.910 1014.260 1796.230 1014.320 ;
        RECT 1795.910 980.460 1796.230 980.520 ;
        RECT 1795.540 980.320 1796.230 980.460 ;
        RECT 1795.540 979.840 1795.680 980.320 ;
        RECT 1795.910 980.260 1796.230 980.320 ;
        RECT 1795.450 979.580 1795.770 979.840 ;
        RECT 1794.530 917.900 1794.850 917.960 ;
        RECT 1795.910 917.900 1796.230 917.960 ;
        RECT 1794.530 917.760 1796.230 917.900 ;
        RECT 1794.530 917.700 1794.850 917.760 ;
        RECT 1795.910 917.700 1796.230 917.760 ;
        RECT 1794.990 869.620 1795.310 869.680 ;
        RECT 1795.910 869.620 1796.230 869.680 ;
        RECT 1794.990 869.480 1796.230 869.620 ;
        RECT 1794.990 869.420 1795.310 869.480 ;
        RECT 1795.910 869.420 1796.230 869.480 ;
        RECT 1794.070 759.120 1794.390 759.180 ;
        RECT 1794.990 759.120 1795.310 759.180 ;
        RECT 1794.070 758.980 1795.310 759.120 ;
        RECT 1794.070 758.920 1794.390 758.980 ;
        RECT 1794.990 758.920 1795.310 758.980 ;
        RECT 1794.070 662.560 1794.390 662.620 ;
        RECT 1794.990 662.560 1795.310 662.620 ;
        RECT 1794.070 662.420 1795.310 662.560 ;
        RECT 1794.070 662.360 1794.390 662.420 ;
        RECT 1794.990 662.360 1795.310 662.420 ;
        RECT 1794.070 566.000 1794.390 566.060 ;
        RECT 1794.990 566.000 1795.310 566.060 ;
        RECT 1794.070 565.860 1795.310 566.000 ;
        RECT 1794.070 565.800 1794.390 565.860 ;
        RECT 1794.990 565.800 1795.310 565.860 ;
        RECT 1794.070 469.440 1794.390 469.500 ;
        RECT 1794.990 469.440 1795.310 469.500 ;
        RECT 1794.070 469.300 1795.310 469.440 ;
        RECT 1794.070 469.240 1794.390 469.300 ;
        RECT 1794.990 469.240 1795.310 469.300 ;
        RECT 1794.070 372.880 1794.390 372.940 ;
        RECT 1794.990 372.880 1795.310 372.940 ;
        RECT 1794.070 372.740 1795.310 372.880 ;
        RECT 1794.070 372.680 1794.390 372.740 ;
        RECT 1794.990 372.680 1795.310 372.740 ;
        RECT 1794.070 276.320 1794.390 276.380 ;
        RECT 1794.990 276.320 1795.310 276.380 ;
        RECT 1794.070 276.180 1795.310 276.320 ;
        RECT 1794.070 276.120 1794.390 276.180 ;
        RECT 1794.990 276.120 1795.310 276.180 ;
        RECT 1794.070 179.760 1794.390 179.820 ;
        RECT 1794.990 179.760 1795.310 179.820 ;
        RECT 1794.070 179.620 1795.310 179.760 ;
        RECT 1794.070 179.560 1794.390 179.620 ;
        RECT 1794.990 179.560 1795.310 179.620 ;
        RECT 1794.070 83.200 1794.390 83.260 ;
        RECT 1794.990 83.200 1795.310 83.260 ;
        RECT 1794.070 83.060 1795.310 83.200 ;
        RECT 1794.070 83.000 1794.390 83.060 ;
        RECT 1794.990 83.000 1795.310 83.060 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 1794.990 17.240 1795.310 17.300 ;
        RECT 2.830 17.100 1795.310 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 1794.990 17.040 1795.310 17.100 ;
      LAYER via ;
        RECT 1796.400 1876.840 1796.660 1877.100 ;
        RECT 1797.780 1876.840 1798.040 1877.100 ;
        RECT 1796.400 1828.220 1796.660 1828.480 ;
        RECT 1795.940 1800.340 1796.200 1800.600 ;
        RECT 1794.100 1676.580 1794.360 1676.840 ;
        RECT 1795.480 1676.580 1795.740 1676.840 ;
        RECT 1794.100 1627.960 1794.360 1628.220 ;
        RECT 1795.480 1627.960 1795.740 1628.220 ;
        RECT 1794.100 1580.020 1794.360 1580.280 ;
        RECT 1795.480 1580.020 1795.740 1580.280 ;
        RECT 1794.100 1531.400 1794.360 1531.660 ;
        RECT 1795.480 1531.400 1795.740 1531.660 ;
        RECT 1794.100 1483.460 1794.360 1483.720 ;
        RECT 1795.480 1483.460 1795.740 1483.720 ;
        RECT 1794.100 1434.840 1794.360 1435.100 ;
        RECT 1795.480 1434.840 1795.740 1435.100 ;
        RECT 1794.100 1386.900 1794.360 1387.160 ;
        RECT 1795.480 1386.900 1795.740 1387.160 ;
        RECT 1794.100 1338.620 1794.360 1338.880 ;
        RECT 1795.020 1338.620 1795.280 1338.880 ;
        RECT 1794.560 1303.940 1794.820 1304.200 ;
        RECT 1794.100 1256.000 1794.360 1256.260 ;
        RECT 1794.560 1207.040 1794.820 1207.300 ;
        RECT 1795.480 1173.040 1795.740 1173.300 ;
        RECT 1794.560 1110.820 1794.820 1111.080 ;
        RECT 1795.940 1110.820 1796.200 1111.080 ;
        RECT 1795.940 1076.820 1796.200 1077.080 ;
        RECT 1795.480 1076.140 1795.740 1076.400 ;
        RECT 1794.560 1014.260 1794.820 1014.520 ;
        RECT 1795.940 1014.260 1796.200 1014.520 ;
        RECT 1795.940 980.260 1796.200 980.520 ;
        RECT 1795.480 979.580 1795.740 979.840 ;
        RECT 1794.560 917.700 1794.820 917.960 ;
        RECT 1795.940 917.700 1796.200 917.960 ;
        RECT 1795.020 869.420 1795.280 869.680 ;
        RECT 1795.940 869.420 1796.200 869.680 ;
        RECT 1794.100 758.920 1794.360 759.180 ;
        RECT 1795.020 758.920 1795.280 759.180 ;
        RECT 1794.100 662.360 1794.360 662.620 ;
        RECT 1795.020 662.360 1795.280 662.620 ;
        RECT 1794.100 565.800 1794.360 566.060 ;
        RECT 1795.020 565.800 1795.280 566.060 ;
        RECT 1794.100 469.240 1794.360 469.500 ;
        RECT 1795.020 469.240 1795.280 469.500 ;
        RECT 1794.100 372.680 1794.360 372.940 ;
        RECT 1795.020 372.680 1795.280 372.940 ;
        RECT 1794.100 276.120 1794.360 276.380 ;
        RECT 1795.020 276.120 1795.280 276.380 ;
        RECT 1794.100 179.560 1794.360 179.820 ;
        RECT 1795.020 179.560 1795.280 179.820 ;
        RECT 1794.100 83.000 1794.360 83.260 ;
        RECT 1795.020 83.000 1795.280 83.260 ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 1795.020 17.040 1795.280 17.300 ;
      LAYER met2 ;
        RECT 1797.770 1877.635 1798.050 1878.005 ;
        RECT 1797.840 1877.130 1797.980 1877.635 ;
        RECT 1796.400 1876.810 1796.660 1877.130 ;
        RECT 1797.780 1876.810 1798.040 1877.130 ;
        RECT 1796.460 1828.510 1796.600 1876.810 ;
        RECT 1796.400 1828.190 1796.660 1828.510 ;
        RECT 1795.940 1800.370 1796.200 1800.630 ;
        RECT 1795.540 1800.310 1796.200 1800.370 ;
        RECT 1795.540 1800.230 1796.140 1800.310 ;
        RECT 1795.540 1676.870 1795.680 1800.230 ;
        RECT 1794.100 1676.550 1794.360 1676.870 ;
        RECT 1795.480 1676.550 1795.740 1676.870 ;
        RECT 1794.160 1628.250 1794.300 1676.550 ;
        RECT 1794.100 1627.930 1794.360 1628.250 ;
        RECT 1795.480 1627.930 1795.740 1628.250 ;
        RECT 1795.540 1580.310 1795.680 1627.930 ;
        RECT 1794.100 1579.990 1794.360 1580.310 ;
        RECT 1795.480 1579.990 1795.740 1580.310 ;
        RECT 1794.160 1531.690 1794.300 1579.990 ;
        RECT 1794.100 1531.370 1794.360 1531.690 ;
        RECT 1795.480 1531.370 1795.740 1531.690 ;
        RECT 1795.540 1483.750 1795.680 1531.370 ;
        RECT 1794.100 1483.430 1794.360 1483.750 ;
        RECT 1795.480 1483.430 1795.740 1483.750 ;
        RECT 1794.160 1435.130 1794.300 1483.430 ;
        RECT 1794.100 1434.810 1794.360 1435.130 ;
        RECT 1795.480 1434.810 1795.740 1435.130 ;
        RECT 1794.160 1387.190 1794.300 1387.345 ;
        RECT 1795.540 1387.190 1795.680 1434.810 ;
        RECT 1794.100 1386.930 1794.360 1387.190 ;
        RECT 1794.100 1386.870 1795.220 1386.930 ;
        RECT 1795.480 1386.870 1795.740 1387.190 ;
        RECT 1794.160 1386.790 1795.220 1386.870 ;
        RECT 1795.080 1338.910 1795.220 1386.790 ;
        RECT 1794.100 1338.650 1794.360 1338.910 ;
        RECT 1794.100 1338.590 1794.760 1338.650 ;
        RECT 1795.020 1338.590 1795.280 1338.910 ;
        RECT 1794.160 1338.510 1794.760 1338.590 ;
        RECT 1794.620 1337.970 1794.760 1338.510 ;
        RECT 1794.620 1337.830 1795.220 1337.970 ;
        RECT 1795.080 1317.570 1795.220 1337.830 ;
        RECT 1794.620 1317.430 1795.220 1317.570 ;
        RECT 1794.620 1304.230 1794.760 1317.430 ;
        RECT 1794.560 1303.910 1794.820 1304.230 ;
        RECT 1794.100 1255.970 1794.360 1256.290 ;
        RECT 1794.160 1221.010 1794.300 1255.970 ;
        RECT 1794.160 1220.870 1794.760 1221.010 ;
        RECT 1794.620 1207.330 1794.760 1220.870 ;
        RECT 1794.560 1207.010 1794.820 1207.330 ;
        RECT 1795.480 1173.010 1795.740 1173.330 ;
        RECT 1795.540 1159.245 1795.680 1173.010 ;
        RECT 1794.550 1158.875 1794.830 1159.245 ;
        RECT 1795.470 1158.875 1795.750 1159.245 ;
        RECT 1794.620 1111.110 1794.760 1158.875 ;
        RECT 1794.560 1110.790 1794.820 1111.110 ;
        RECT 1795.940 1110.790 1796.200 1111.110 ;
        RECT 1796.000 1077.110 1796.140 1110.790 ;
        RECT 1795.940 1076.790 1796.200 1077.110 ;
        RECT 1795.480 1076.110 1795.740 1076.430 ;
        RECT 1795.540 1062.685 1795.680 1076.110 ;
        RECT 1794.550 1062.315 1794.830 1062.685 ;
        RECT 1795.470 1062.315 1795.750 1062.685 ;
        RECT 1794.620 1014.550 1794.760 1062.315 ;
        RECT 1794.560 1014.230 1794.820 1014.550 ;
        RECT 1795.940 1014.230 1796.200 1014.550 ;
        RECT 1796.000 980.550 1796.140 1014.230 ;
        RECT 1795.940 980.230 1796.200 980.550 ;
        RECT 1795.480 979.550 1795.740 979.870 ;
        RECT 1795.540 966.125 1795.680 979.550 ;
        RECT 1794.550 965.755 1794.830 966.125 ;
        RECT 1795.470 965.755 1795.750 966.125 ;
        RECT 1794.620 917.990 1794.760 965.755 ;
        RECT 1794.560 917.670 1794.820 917.990 ;
        RECT 1795.940 917.670 1796.200 917.990 ;
        RECT 1796.000 869.710 1796.140 917.670 ;
        RECT 1795.020 869.565 1795.280 869.710 ;
        RECT 1793.630 869.195 1793.910 869.565 ;
        RECT 1795.010 869.195 1795.290 869.565 ;
        RECT 1795.940 869.390 1796.200 869.710 ;
        RECT 1793.700 821.285 1793.840 869.195 ;
        RECT 1793.630 820.915 1793.910 821.285 ;
        RECT 1794.550 820.915 1794.830 821.285 ;
        RECT 1794.620 807.570 1794.760 820.915 ;
        RECT 1794.620 807.430 1795.220 807.570 ;
        RECT 1795.080 759.210 1795.220 807.430 ;
        RECT 1794.100 758.890 1794.360 759.210 ;
        RECT 1795.020 758.890 1795.280 759.210 ;
        RECT 1794.160 758.610 1794.300 758.890 ;
        RECT 1794.160 758.470 1794.760 758.610 ;
        RECT 1794.620 711.010 1794.760 758.470 ;
        RECT 1794.620 710.870 1795.220 711.010 ;
        RECT 1795.080 662.650 1795.220 710.870 ;
        RECT 1794.100 662.330 1794.360 662.650 ;
        RECT 1795.020 662.330 1795.280 662.650 ;
        RECT 1794.160 662.050 1794.300 662.330 ;
        RECT 1794.160 661.910 1794.760 662.050 ;
        RECT 1794.620 614.450 1794.760 661.910 ;
        RECT 1794.620 614.310 1795.220 614.450 ;
        RECT 1795.080 566.090 1795.220 614.310 ;
        RECT 1794.100 565.770 1794.360 566.090 ;
        RECT 1795.020 565.770 1795.280 566.090 ;
        RECT 1794.160 565.490 1794.300 565.770 ;
        RECT 1794.160 565.350 1794.760 565.490 ;
        RECT 1794.620 517.890 1794.760 565.350 ;
        RECT 1794.620 517.750 1795.220 517.890 ;
        RECT 1795.080 469.530 1795.220 517.750 ;
        RECT 1794.100 469.210 1794.360 469.530 ;
        RECT 1795.020 469.210 1795.280 469.530 ;
        RECT 1794.160 468.930 1794.300 469.210 ;
        RECT 1794.160 468.790 1794.760 468.930 ;
        RECT 1794.620 421.330 1794.760 468.790 ;
        RECT 1794.620 421.190 1795.220 421.330 ;
        RECT 1795.080 372.970 1795.220 421.190 ;
        RECT 1794.100 372.650 1794.360 372.970 ;
        RECT 1795.020 372.650 1795.280 372.970 ;
        RECT 1794.160 372.370 1794.300 372.650 ;
        RECT 1794.160 372.230 1794.760 372.370 ;
        RECT 1794.620 324.770 1794.760 372.230 ;
        RECT 1794.620 324.630 1795.220 324.770 ;
        RECT 1795.080 276.410 1795.220 324.630 ;
        RECT 1794.100 276.090 1794.360 276.410 ;
        RECT 1795.020 276.090 1795.280 276.410 ;
        RECT 1794.160 275.810 1794.300 276.090 ;
        RECT 1794.160 275.670 1794.760 275.810 ;
        RECT 1794.620 228.210 1794.760 275.670 ;
        RECT 1794.620 228.070 1795.220 228.210 ;
        RECT 1795.080 179.850 1795.220 228.070 ;
        RECT 1794.100 179.530 1794.360 179.850 ;
        RECT 1795.020 179.530 1795.280 179.850 ;
        RECT 1794.160 130.970 1794.300 179.530 ;
        RECT 1794.160 130.830 1795.220 130.970 ;
        RECT 1795.080 83.290 1795.220 130.830 ;
        RECT 1794.100 82.970 1794.360 83.290 ;
        RECT 1795.020 82.970 1795.280 83.290 ;
        RECT 1794.160 34.410 1794.300 82.970 ;
        RECT 1794.160 34.270 1795.220 34.410 ;
        RECT 1795.080 17.330 1795.220 34.270 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 1795.020 17.010 1795.280 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 1797.770 1877.680 1798.050 1877.960 ;
        RECT 1794.550 1158.920 1794.830 1159.200 ;
        RECT 1795.470 1158.920 1795.750 1159.200 ;
        RECT 1794.550 1062.360 1794.830 1062.640 ;
        RECT 1795.470 1062.360 1795.750 1062.640 ;
        RECT 1794.550 965.800 1794.830 966.080 ;
        RECT 1795.470 965.800 1795.750 966.080 ;
        RECT 1793.630 869.240 1793.910 869.520 ;
        RECT 1795.010 869.240 1795.290 869.520 ;
        RECT 1793.630 820.960 1793.910 821.240 ;
        RECT 1794.550 820.960 1794.830 821.240 ;
      LAYER met3 ;
        RECT 1797.000 1880.240 1801.000 1880.840 ;
        RECT 1797.990 1877.985 1798.290 1880.240 ;
        RECT 1797.745 1877.670 1798.290 1877.985 ;
        RECT 1797.745 1877.655 1798.075 1877.670 ;
        RECT 1794.525 1159.210 1794.855 1159.225 ;
        RECT 1795.445 1159.210 1795.775 1159.225 ;
        RECT 1794.525 1158.910 1795.775 1159.210 ;
        RECT 1794.525 1158.895 1794.855 1158.910 ;
        RECT 1795.445 1158.895 1795.775 1158.910 ;
        RECT 1794.525 1062.650 1794.855 1062.665 ;
        RECT 1795.445 1062.650 1795.775 1062.665 ;
        RECT 1794.525 1062.350 1795.775 1062.650 ;
        RECT 1794.525 1062.335 1794.855 1062.350 ;
        RECT 1795.445 1062.335 1795.775 1062.350 ;
        RECT 1794.525 966.090 1794.855 966.105 ;
        RECT 1795.445 966.090 1795.775 966.105 ;
        RECT 1794.525 965.790 1795.775 966.090 ;
        RECT 1794.525 965.775 1794.855 965.790 ;
        RECT 1795.445 965.775 1795.775 965.790 ;
        RECT 1793.605 869.530 1793.935 869.545 ;
        RECT 1794.985 869.530 1795.315 869.545 ;
        RECT 1793.605 869.230 1795.315 869.530 ;
        RECT 1793.605 869.215 1793.935 869.230 ;
        RECT 1794.985 869.215 1795.315 869.230 ;
        RECT 1793.605 821.250 1793.935 821.265 ;
        RECT 1794.525 821.250 1794.855 821.265 ;
        RECT 1793.605 820.950 1794.855 821.250 ;
        RECT 1793.605 820.935 1793.935 820.950 ;
        RECT 1794.525 820.935 1794.855 820.950 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.930 -4.570 -7.030 3524.250 ;
        RECT 4.070 -9.170 6.970 3528.850 ;
        RECT 184.070 -9.170 186.970 3528.850 ;
        RECT 364.070 -9.170 366.970 3528.850 ;
        RECT 544.070 -9.170 546.970 3528.850 ;
        RECT 724.070 -9.170 726.970 3528.850 ;
        RECT 904.070 -9.170 906.970 3528.850 ;
        RECT 1084.070 -9.170 1086.970 3528.850 ;
        RECT 1264.070 -9.170 1266.970 3528.850 ;
        RECT 1444.070 -9.170 1446.970 3528.850 ;
        RECT 1624.070 -9.170 1626.970 3528.850 ;
        RECT 1804.070 -9.170 1806.970 3528.850 ;
        RECT 1984.070 -9.170 1986.970 3528.850 ;
        RECT 2164.070 -9.170 2166.970 3528.850 ;
        RECT 2344.070 -9.170 2346.970 3528.850 ;
        RECT 2524.070 -9.170 2526.970 3528.850 ;
        RECT 2704.070 -9.170 2706.970 3528.850 ;
        RECT 2884.070 -9.170 2886.970 3528.850 ;
        RECT 2926.650 -4.570 2929.550 3524.250 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.930 3524.250 -7.030 3524.310 ;
        RECT 4.070 3524.250 6.970 3524.310 ;
        RECT 184.070 3524.250 186.970 3524.310 ;
        RECT 364.070 3524.250 366.970 3524.310 ;
        RECT 544.070 3524.250 546.970 3524.310 ;
        RECT 724.070 3524.250 726.970 3524.310 ;
        RECT 904.070 3524.250 906.970 3524.310 ;
        RECT 1084.070 3524.250 1086.970 3524.310 ;
        RECT 1264.070 3524.250 1266.970 3524.310 ;
        RECT 1444.070 3524.250 1446.970 3524.310 ;
        RECT 1624.070 3524.250 1626.970 3524.310 ;
        RECT 1804.070 3524.250 1806.970 3524.310 ;
        RECT 1984.070 3524.250 1986.970 3524.310 ;
        RECT 2164.070 3524.250 2166.970 3524.310 ;
        RECT 2344.070 3524.250 2346.970 3524.310 ;
        RECT 2524.070 3524.250 2526.970 3524.310 ;
        RECT 2704.070 3524.250 2706.970 3524.310 ;
        RECT 2884.070 3524.250 2886.970 3524.310 ;
        RECT 2926.650 3524.250 2929.550 3524.310 ;
        RECT -9.930 3521.350 2929.550 3524.250 ;
        RECT -9.930 3521.290 -7.030 3521.350 ;
        RECT 4.070 3521.290 6.970 3521.350 ;
        RECT 184.070 3521.290 186.970 3521.350 ;
        RECT 364.070 3521.290 366.970 3521.350 ;
        RECT 544.070 3521.290 546.970 3521.350 ;
        RECT 724.070 3521.290 726.970 3521.350 ;
        RECT 904.070 3521.290 906.970 3521.350 ;
        RECT 1084.070 3521.290 1086.970 3521.350 ;
        RECT 1264.070 3521.290 1266.970 3521.350 ;
        RECT 1444.070 3521.290 1446.970 3521.350 ;
        RECT 1624.070 3521.290 1626.970 3521.350 ;
        RECT 1804.070 3521.290 1806.970 3521.350 ;
        RECT 1984.070 3521.290 1986.970 3521.350 ;
        RECT 2164.070 3521.290 2166.970 3521.350 ;
        RECT 2344.070 3521.290 2346.970 3521.350 ;
        RECT 2524.070 3521.290 2526.970 3521.350 ;
        RECT 2704.070 3521.290 2706.970 3521.350 ;
        RECT 2884.070 3521.290 2886.970 3521.350 ;
        RECT 2926.650 3521.290 2929.550 3521.350 ;
        RECT -9.930 3432.330 -7.030 3432.390 ;
        RECT 4.070 3432.330 6.970 3432.390 ;
        RECT 184.070 3432.330 186.970 3432.390 ;
        RECT 364.070 3432.330 366.970 3432.390 ;
        RECT 544.070 3432.330 546.970 3432.390 ;
        RECT 724.070 3432.330 726.970 3432.390 ;
        RECT 904.070 3432.330 906.970 3432.390 ;
        RECT 1084.070 3432.330 1086.970 3432.390 ;
        RECT 1264.070 3432.330 1266.970 3432.390 ;
        RECT 1444.070 3432.330 1446.970 3432.390 ;
        RECT 1624.070 3432.330 1626.970 3432.390 ;
        RECT 1804.070 3432.330 1806.970 3432.390 ;
        RECT 1984.070 3432.330 1986.970 3432.390 ;
        RECT 2164.070 3432.330 2166.970 3432.390 ;
        RECT 2344.070 3432.330 2346.970 3432.390 ;
        RECT 2524.070 3432.330 2526.970 3432.390 ;
        RECT 2704.070 3432.330 2706.970 3432.390 ;
        RECT 2884.070 3432.330 2886.970 3432.390 ;
        RECT 2926.650 3432.330 2929.550 3432.390 ;
        RECT -14.530 3429.430 2934.150 3432.330 ;
        RECT -9.930 3429.370 -7.030 3429.430 ;
        RECT 4.070 3429.370 6.970 3429.430 ;
        RECT 184.070 3429.370 186.970 3429.430 ;
        RECT 364.070 3429.370 366.970 3429.430 ;
        RECT 544.070 3429.370 546.970 3429.430 ;
        RECT 724.070 3429.370 726.970 3429.430 ;
        RECT 904.070 3429.370 906.970 3429.430 ;
        RECT 1084.070 3429.370 1086.970 3429.430 ;
        RECT 1264.070 3429.370 1266.970 3429.430 ;
        RECT 1444.070 3429.370 1446.970 3429.430 ;
        RECT 1624.070 3429.370 1626.970 3429.430 ;
        RECT 1804.070 3429.370 1806.970 3429.430 ;
        RECT 1984.070 3429.370 1986.970 3429.430 ;
        RECT 2164.070 3429.370 2166.970 3429.430 ;
        RECT 2344.070 3429.370 2346.970 3429.430 ;
        RECT 2524.070 3429.370 2526.970 3429.430 ;
        RECT 2704.070 3429.370 2706.970 3429.430 ;
        RECT 2884.070 3429.370 2886.970 3429.430 ;
        RECT 2926.650 3429.370 2929.550 3429.430 ;
        RECT -9.930 3252.330 -7.030 3252.390 ;
        RECT 4.070 3252.330 6.970 3252.390 ;
        RECT 184.070 3252.330 186.970 3252.390 ;
        RECT 364.070 3252.330 366.970 3252.390 ;
        RECT 544.070 3252.330 546.970 3252.390 ;
        RECT 724.070 3252.330 726.970 3252.390 ;
        RECT 904.070 3252.330 906.970 3252.390 ;
        RECT 1084.070 3252.330 1086.970 3252.390 ;
        RECT 1264.070 3252.330 1266.970 3252.390 ;
        RECT 1444.070 3252.330 1446.970 3252.390 ;
        RECT 1624.070 3252.330 1626.970 3252.390 ;
        RECT 1804.070 3252.330 1806.970 3252.390 ;
        RECT 1984.070 3252.330 1986.970 3252.390 ;
        RECT 2164.070 3252.330 2166.970 3252.390 ;
        RECT 2344.070 3252.330 2346.970 3252.390 ;
        RECT 2524.070 3252.330 2526.970 3252.390 ;
        RECT 2704.070 3252.330 2706.970 3252.390 ;
        RECT 2884.070 3252.330 2886.970 3252.390 ;
        RECT 2926.650 3252.330 2929.550 3252.390 ;
        RECT -14.530 3249.430 2934.150 3252.330 ;
        RECT -9.930 3249.370 -7.030 3249.430 ;
        RECT 4.070 3249.370 6.970 3249.430 ;
        RECT 184.070 3249.370 186.970 3249.430 ;
        RECT 364.070 3249.370 366.970 3249.430 ;
        RECT 544.070 3249.370 546.970 3249.430 ;
        RECT 724.070 3249.370 726.970 3249.430 ;
        RECT 904.070 3249.370 906.970 3249.430 ;
        RECT 1084.070 3249.370 1086.970 3249.430 ;
        RECT 1264.070 3249.370 1266.970 3249.430 ;
        RECT 1444.070 3249.370 1446.970 3249.430 ;
        RECT 1624.070 3249.370 1626.970 3249.430 ;
        RECT 1804.070 3249.370 1806.970 3249.430 ;
        RECT 1984.070 3249.370 1986.970 3249.430 ;
        RECT 2164.070 3249.370 2166.970 3249.430 ;
        RECT 2344.070 3249.370 2346.970 3249.430 ;
        RECT 2524.070 3249.370 2526.970 3249.430 ;
        RECT 2704.070 3249.370 2706.970 3249.430 ;
        RECT 2884.070 3249.370 2886.970 3249.430 ;
        RECT 2926.650 3249.370 2929.550 3249.430 ;
        RECT -9.930 3072.330 -7.030 3072.390 ;
        RECT 4.070 3072.330 6.970 3072.390 ;
        RECT 184.070 3072.330 186.970 3072.390 ;
        RECT 364.070 3072.330 366.970 3072.390 ;
        RECT 544.070 3072.330 546.970 3072.390 ;
        RECT 724.070 3072.330 726.970 3072.390 ;
        RECT 904.070 3072.330 906.970 3072.390 ;
        RECT 1084.070 3072.330 1086.970 3072.390 ;
        RECT 1264.070 3072.330 1266.970 3072.390 ;
        RECT 1444.070 3072.330 1446.970 3072.390 ;
        RECT 1624.070 3072.330 1626.970 3072.390 ;
        RECT 1804.070 3072.330 1806.970 3072.390 ;
        RECT 1984.070 3072.330 1986.970 3072.390 ;
        RECT 2164.070 3072.330 2166.970 3072.390 ;
        RECT 2344.070 3072.330 2346.970 3072.390 ;
        RECT 2524.070 3072.330 2526.970 3072.390 ;
        RECT 2704.070 3072.330 2706.970 3072.390 ;
        RECT 2884.070 3072.330 2886.970 3072.390 ;
        RECT 2926.650 3072.330 2929.550 3072.390 ;
        RECT -14.530 3069.430 2934.150 3072.330 ;
        RECT -9.930 3069.370 -7.030 3069.430 ;
        RECT 4.070 3069.370 6.970 3069.430 ;
        RECT 184.070 3069.370 186.970 3069.430 ;
        RECT 364.070 3069.370 366.970 3069.430 ;
        RECT 544.070 3069.370 546.970 3069.430 ;
        RECT 724.070 3069.370 726.970 3069.430 ;
        RECT 904.070 3069.370 906.970 3069.430 ;
        RECT 1084.070 3069.370 1086.970 3069.430 ;
        RECT 1264.070 3069.370 1266.970 3069.430 ;
        RECT 1444.070 3069.370 1446.970 3069.430 ;
        RECT 1624.070 3069.370 1626.970 3069.430 ;
        RECT 1804.070 3069.370 1806.970 3069.430 ;
        RECT 1984.070 3069.370 1986.970 3069.430 ;
        RECT 2164.070 3069.370 2166.970 3069.430 ;
        RECT 2344.070 3069.370 2346.970 3069.430 ;
        RECT 2524.070 3069.370 2526.970 3069.430 ;
        RECT 2704.070 3069.370 2706.970 3069.430 ;
        RECT 2884.070 3069.370 2886.970 3069.430 ;
        RECT 2926.650 3069.370 2929.550 3069.430 ;
        RECT -9.930 2892.330 -7.030 2892.390 ;
        RECT 4.070 2892.330 6.970 2892.390 ;
        RECT 184.070 2892.330 186.970 2892.390 ;
        RECT 364.070 2892.330 366.970 2892.390 ;
        RECT 544.070 2892.330 546.970 2892.390 ;
        RECT 724.070 2892.330 726.970 2892.390 ;
        RECT 904.070 2892.330 906.970 2892.390 ;
        RECT 1084.070 2892.330 1086.970 2892.390 ;
        RECT 1264.070 2892.330 1266.970 2892.390 ;
        RECT 1444.070 2892.330 1446.970 2892.390 ;
        RECT 1624.070 2892.330 1626.970 2892.390 ;
        RECT 1804.070 2892.330 1806.970 2892.390 ;
        RECT 1984.070 2892.330 1986.970 2892.390 ;
        RECT 2164.070 2892.330 2166.970 2892.390 ;
        RECT 2344.070 2892.330 2346.970 2892.390 ;
        RECT 2524.070 2892.330 2526.970 2892.390 ;
        RECT 2704.070 2892.330 2706.970 2892.390 ;
        RECT 2884.070 2892.330 2886.970 2892.390 ;
        RECT 2926.650 2892.330 2929.550 2892.390 ;
        RECT -14.530 2889.430 2934.150 2892.330 ;
        RECT -9.930 2889.370 -7.030 2889.430 ;
        RECT 4.070 2889.370 6.970 2889.430 ;
        RECT 184.070 2889.370 186.970 2889.430 ;
        RECT 364.070 2889.370 366.970 2889.430 ;
        RECT 544.070 2889.370 546.970 2889.430 ;
        RECT 724.070 2889.370 726.970 2889.430 ;
        RECT 904.070 2889.370 906.970 2889.430 ;
        RECT 1084.070 2889.370 1086.970 2889.430 ;
        RECT 1264.070 2889.370 1266.970 2889.430 ;
        RECT 1444.070 2889.370 1446.970 2889.430 ;
        RECT 1624.070 2889.370 1626.970 2889.430 ;
        RECT 1804.070 2889.370 1806.970 2889.430 ;
        RECT 1984.070 2889.370 1986.970 2889.430 ;
        RECT 2164.070 2889.370 2166.970 2889.430 ;
        RECT 2344.070 2889.370 2346.970 2889.430 ;
        RECT 2524.070 2889.370 2526.970 2889.430 ;
        RECT 2704.070 2889.370 2706.970 2889.430 ;
        RECT 2884.070 2889.370 2886.970 2889.430 ;
        RECT 2926.650 2889.370 2929.550 2889.430 ;
        RECT -9.930 2712.330 -7.030 2712.390 ;
        RECT 4.070 2712.330 6.970 2712.390 ;
        RECT 184.070 2712.330 186.970 2712.390 ;
        RECT 364.070 2712.330 366.970 2712.390 ;
        RECT 544.070 2712.330 546.970 2712.390 ;
        RECT 724.070 2712.330 726.970 2712.390 ;
        RECT 904.070 2712.330 906.970 2712.390 ;
        RECT 1084.070 2712.330 1086.970 2712.390 ;
        RECT 1264.070 2712.330 1266.970 2712.390 ;
        RECT 1444.070 2712.330 1446.970 2712.390 ;
        RECT 1624.070 2712.330 1626.970 2712.390 ;
        RECT 1804.070 2712.330 1806.970 2712.390 ;
        RECT 1984.070 2712.330 1986.970 2712.390 ;
        RECT 2164.070 2712.330 2166.970 2712.390 ;
        RECT 2344.070 2712.330 2346.970 2712.390 ;
        RECT 2524.070 2712.330 2526.970 2712.390 ;
        RECT 2704.070 2712.330 2706.970 2712.390 ;
        RECT 2884.070 2712.330 2886.970 2712.390 ;
        RECT 2926.650 2712.330 2929.550 2712.390 ;
        RECT -14.530 2709.430 2934.150 2712.330 ;
        RECT -9.930 2709.370 -7.030 2709.430 ;
        RECT 4.070 2709.370 6.970 2709.430 ;
        RECT 184.070 2709.370 186.970 2709.430 ;
        RECT 364.070 2709.370 366.970 2709.430 ;
        RECT 544.070 2709.370 546.970 2709.430 ;
        RECT 724.070 2709.370 726.970 2709.430 ;
        RECT 904.070 2709.370 906.970 2709.430 ;
        RECT 1084.070 2709.370 1086.970 2709.430 ;
        RECT 1264.070 2709.370 1266.970 2709.430 ;
        RECT 1444.070 2709.370 1446.970 2709.430 ;
        RECT 1624.070 2709.370 1626.970 2709.430 ;
        RECT 1804.070 2709.370 1806.970 2709.430 ;
        RECT 1984.070 2709.370 1986.970 2709.430 ;
        RECT 2164.070 2709.370 2166.970 2709.430 ;
        RECT 2344.070 2709.370 2346.970 2709.430 ;
        RECT 2524.070 2709.370 2526.970 2709.430 ;
        RECT 2704.070 2709.370 2706.970 2709.430 ;
        RECT 2884.070 2709.370 2886.970 2709.430 ;
        RECT 2926.650 2709.370 2929.550 2709.430 ;
        RECT -9.930 2532.330 -7.030 2532.390 ;
        RECT 4.070 2532.330 6.970 2532.390 ;
        RECT 184.070 2532.330 186.970 2532.390 ;
        RECT 364.070 2532.330 366.970 2532.390 ;
        RECT 544.070 2532.330 546.970 2532.390 ;
        RECT 724.070 2532.330 726.970 2532.390 ;
        RECT 904.070 2532.330 906.970 2532.390 ;
        RECT 1084.070 2532.330 1086.970 2532.390 ;
        RECT 1264.070 2532.330 1266.970 2532.390 ;
        RECT 1444.070 2532.330 1446.970 2532.390 ;
        RECT 1624.070 2532.330 1626.970 2532.390 ;
        RECT 1804.070 2532.330 1806.970 2532.390 ;
        RECT 1984.070 2532.330 1986.970 2532.390 ;
        RECT 2164.070 2532.330 2166.970 2532.390 ;
        RECT 2344.070 2532.330 2346.970 2532.390 ;
        RECT 2524.070 2532.330 2526.970 2532.390 ;
        RECT 2704.070 2532.330 2706.970 2532.390 ;
        RECT 2884.070 2532.330 2886.970 2532.390 ;
        RECT 2926.650 2532.330 2929.550 2532.390 ;
        RECT -14.530 2529.430 2934.150 2532.330 ;
        RECT -9.930 2529.370 -7.030 2529.430 ;
        RECT 4.070 2529.370 6.970 2529.430 ;
        RECT 184.070 2529.370 186.970 2529.430 ;
        RECT 364.070 2529.370 366.970 2529.430 ;
        RECT 544.070 2529.370 546.970 2529.430 ;
        RECT 724.070 2529.370 726.970 2529.430 ;
        RECT 904.070 2529.370 906.970 2529.430 ;
        RECT 1084.070 2529.370 1086.970 2529.430 ;
        RECT 1264.070 2529.370 1266.970 2529.430 ;
        RECT 1444.070 2529.370 1446.970 2529.430 ;
        RECT 1624.070 2529.370 1626.970 2529.430 ;
        RECT 1804.070 2529.370 1806.970 2529.430 ;
        RECT 1984.070 2529.370 1986.970 2529.430 ;
        RECT 2164.070 2529.370 2166.970 2529.430 ;
        RECT 2344.070 2529.370 2346.970 2529.430 ;
        RECT 2524.070 2529.370 2526.970 2529.430 ;
        RECT 2704.070 2529.370 2706.970 2529.430 ;
        RECT 2884.070 2529.370 2886.970 2529.430 ;
        RECT 2926.650 2529.370 2929.550 2529.430 ;
        RECT -9.930 2352.330 -7.030 2352.390 ;
        RECT 4.070 2352.330 6.970 2352.390 ;
        RECT 184.070 2352.330 186.970 2352.390 ;
        RECT 364.070 2352.330 366.970 2352.390 ;
        RECT 544.070 2352.330 546.970 2352.390 ;
        RECT 724.070 2352.330 726.970 2352.390 ;
        RECT 904.070 2352.330 906.970 2352.390 ;
        RECT 1084.070 2352.330 1086.970 2352.390 ;
        RECT 1264.070 2352.330 1266.970 2352.390 ;
        RECT 1444.070 2352.330 1446.970 2352.390 ;
        RECT 1624.070 2352.330 1626.970 2352.390 ;
        RECT 1804.070 2352.330 1806.970 2352.390 ;
        RECT 1984.070 2352.330 1986.970 2352.390 ;
        RECT 2164.070 2352.330 2166.970 2352.390 ;
        RECT 2344.070 2352.330 2346.970 2352.390 ;
        RECT 2524.070 2352.330 2526.970 2352.390 ;
        RECT 2704.070 2352.330 2706.970 2352.390 ;
        RECT 2884.070 2352.330 2886.970 2352.390 ;
        RECT 2926.650 2352.330 2929.550 2352.390 ;
        RECT -14.530 2349.430 2934.150 2352.330 ;
        RECT -9.930 2349.370 -7.030 2349.430 ;
        RECT 4.070 2349.370 6.970 2349.430 ;
        RECT 184.070 2349.370 186.970 2349.430 ;
        RECT 364.070 2349.370 366.970 2349.430 ;
        RECT 544.070 2349.370 546.970 2349.430 ;
        RECT 724.070 2349.370 726.970 2349.430 ;
        RECT 904.070 2349.370 906.970 2349.430 ;
        RECT 1084.070 2349.370 1086.970 2349.430 ;
        RECT 1264.070 2349.370 1266.970 2349.430 ;
        RECT 1444.070 2349.370 1446.970 2349.430 ;
        RECT 1624.070 2349.370 1626.970 2349.430 ;
        RECT 1804.070 2349.370 1806.970 2349.430 ;
        RECT 1984.070 2349.370 1986.970 2349.430 ;
        RECT 2164.070 2349.370 2166.970 2349.430 ;
        RECT 2344.070 2349.370 2346.970 2349.430 ;
        RECT 2524.070 2349.370 2526.970 2349.430 ;
        RECT 2704.070 2349.370 2706.970 2349.430 ;
        RECT 2884.070 2349.370 2886.970 2349.430 ;
        RECT 2926.650 2349.370 2929.550 2349.430 ;
        RECT -9.930 2172.330 -7.030 2172.390 ;
        RECT 4.070 2172.330 6.970 2172.390 ;
        RECT 184.070 2172.330 186.970 2172.390 ;
        RECT 364.070 2172.330 366.970 2172.390 ;
        RECT 544.070 2172.330 546.970 2172.390 ;
        RECT 724.070 2172.330 726.970 2172.390 ;
        RECT 904.070 2172.330 906.970 2172.390 ;
        RECT 1084.070 2172.330 1086.970 2172.390 ;
        RECT 1264.070 2172.330 1266.970 2172.390 ;
        RECT 1444.070 2172.330 1446.970 2172.390 ;
        RECT 1624.070 2172.330 1626.970 2172.390 ;
        RECT 1804.070 2172.330 1806.970 2172.390 ;
        RECT 1984.070 2172.330 1986.970 2172.390 ;
        RECT 2164.070 2172.330 2166.970 2172.390 ;
        RECT 2344.070 2172.330 2346.970 2172.390 ;
        RECT 2524.070 2172.330 2526.970 2172.390 ;
        RECT 2704.070 2172.330 2706.970 2172.390 ;
        RECT 2884.070 2172.330 2886.970 2172.390 ;
        RECT 2926.650 2172.330 2929.550 2172.390 ;
        RECT -14.530 2169.430 2934.150 2172.330 ;
        RECT -9.930 2169.370 -7.030 2169.430 ;
        RECT 4.070 2169.370 6.970 2169.430 ;
        RECT 184.070 2169.370 186.970 2169.430 ;
        RECT 364.070 2169.370 366.970 2169.430 ;
        RECT 544.070 2169.370 546.970 2169.430 ;
        RECT 724.070 2169.370 726.970 2169.430 ;
        RECT 904.070 2169.370 906.970 2169.430 ;
        RECT 1084.070 2169.370 1086.970 2169.430 ;
        RECT 1264.070 2169.370 1266.970 2169.430 ;
        RECT 1444.070 2169.370 1446.970 2169.430 ;
        RECT 1624.070 2169.370 1626.970 2169.430 ;
        RECT 1804.070 2169.370 1806.970 2169.430 ;
        RECT 1984.070 2169.370 1986.970 2169.430 ;
        RECT 2164.070 2169.370 2166.970 2169.430 ;
        RECT 2344.070 2169.370 2346.970 2169.430 ;
        RECT 2524.070 2169.370 2526.970 2169.430 ;
        RECT 2704.070 2169.370 2706.970 2169.430 ;
        RECT 2884.070 2169.370 2886.970 2169.430 ;
        RECT 2926.650 2169.370 2929.550 2169.430 ;
        RECT -9.930 1992.330 -7.030 1992.390 ;
        RECT 4.070 1992.330 6.970 1992.390 ;
        RECT 184.070 1992.330 186.970 1992.390 ;
        RECT 364.070 1992.330 366.970 1992.390 ;
        RECT 544.070 1992.330 546.970 1992.390 ;
        RECT 724.070 1992.330 726.970 1992.390 ;
        RECT 904.070 1992.330 906.970 1992.390 ;
        RECT 1084.070 1992.330 1086.970 1992.390 ;
        RECT 1264.070 1992.330 1266.970 1992.390 ;
        RECT 1444.070 1992.330 1446.970 1992.390 ;
        RECT 1624.070 1992.330 1626.970 1992.390 ;
        RECT 1804.070 1992.330 1806.970 1992.390 ;
        RECT 1984.070 1992.330 1986.970 1992.390 ;
        RECT 2164.070 1992.330 2166.970 1992.390 ;
        RECT 2344.070 1992.330 2346.970 1992.390 ;
        RECT 2524.070 1992.330 2526.970 1992.390 ;
        RECT 2704.070 1992.330 2706.970 1992.390 ;
        RECT 2884.070 1992.330 2886.970 1992.390 ;
        RECT 2926.650 1992.330 2929.550 1992.390 ;
        RECT -14.530 1989.430 2934.150 1992.330 ;
        RECT -9.930 1989.370 -7.030 1989.430 ;
        RECT 4.070 1989.370 6.970 1989.430 ;
        RECT 184.070 1989.370 186.970 1989.430 ;
        RECT 364.070 1989.370 366.970 1989.430 ;
        RECT 544.070 1989.370 546.970 1989.430 ;
        RECT 724.070 1989.370 726.970 1989.430 ;
        RECT 904.070 1989.370 906.970 1989.430 ;
        RECT 1084.070 1989.370 1086.970 1989.430 ;
        RECT 1264.070 1989.370 1266.970 1989.430 ;
        RECT 1444.070 1989.370 1446.970 1989.430 ;
        RECT 1624.070 1989.370 1626.970 1989.430 ;
        RECT 1804.070 1989.370 1806.970 1989.430 ;
        RECT 1984.070 1989.370 1986.970 1989.430 ;
        RECT 2164.070 1989.370 2166.970 1989.430 ;
        RECT 2344.070 1989.370 2346.970 1989.430 ;
        RECT 2524.070 1989.370 2526.970 1989.430 ;
        RECT 2704.070 1989.370 2706.970 1989.430 ;
        RECT 2884.070 1989.370 2886.970 1989.430 ;
        RECT 2926.650 1989.370 2929.550 1989.430 ;
        RECT -9.930 1812.330 -7.030 1812.390 ;
        RECT 4.070 1812.330 6.970 1812.390 ;
        RECT 184.070 1812.330 186.970 1812.390 ;
        RECT 364.070 1812.330 366.970 1812.390 ;
        RECT 544.070 1812.330 546.970 1812.390 ;
        RECT 724.070 1812.330 726.970 1812.390 ;
        RECT 904.070 1812.330 906.970 1812.390 ;
        RECT 1084.070 1812.330 1086.970 1812.390 ;
        RECT 1264.070 1812.330 1266.970 1812.390 ;
        RECT 1444.070 1812.330 1446.970 1812.390 ;
        RECT 1624.070 1812.330 1626.970 1812.390 ;
        RECT 1804.070 1812.330 1806.970 1812.390 ;
        RECT 1984.070 1812.330 1986.970 1812.390 ;
        RECT 2164.070 1812.330 2166.970 1812.390 ;
        RECT 2344.070 1812.330 2346.970 1812.390 ;
        RECT 2524.070 1812.330 2526.970 1812.390 ;
        RECT 2704.070 1812.330 2706.970 1812.390 ;
        RECT 2884.070 1812.330 2886.970 1812.390 ;
        RECT 2926.650 1812.330 2929.550 1812.390 ;
        RECT -14.530 1809.430 2934.150 1812.330 ;
        RECT -9.930 1809.370 -7.030 1809.430 ;
        RECT 4.070 1809.370 6.970 1809.430 ;
        RECT 184.070 1809.370 186.970 1809.430 ;
        RECT 364.070 1809.370 366.970 1809.430 ;
        RECT 544.070 1809.370 546.970 1809.430 ;
        RECT 724.070 1809.370 726.970 1809.430 ;
        RECT 904.070 1809.370 906.970 1809.430 ;
        RECT 1084.070 1809.370 1086.970 1809.430 ;
        RECT 1264.070 1809.370 1266.970 1809.430 ;
        RECT 1444.070 1809.370 1446.970 1809.430 ;
        RECT 1624.070 1809.370 1626.970 1809.430 ;
        RECT 1804.070 1809.370 1806.970 1809.430 ;
        RECT 1984.070 1809.370 1986.970 1809.430 ;
        RECT 2164.070 1809.370 2166.970 1809.430 ;
        RECT 2344.070 1809.370 2346.970 1809.430 ;
        RECT 2524.070 1809.370 2526.970 1809.430 ;
        RECT 2704.070 1809.370 2706.970 1809.430 ;
        RECT 2884.070 1809.370 2886.970 1809.430 ;
        RECT 2926.650 1809.370 2929.550 1809.430 ;
        RECT -9.930 1632.330 -7.030 1632.390 ;
        RECT 4.070 1632.330 6.970 1632.390 ;
        RECT 184.070 1632.330 186.970 1632.390 ;
        RECT 364.070 1632.330 366.970 1632.390 ;
        RECT 544.070 1632.330 546.970 1632.390 ;
        RECT 724.070 1632.330 726.970 1632.390 ;
        RECT 904.070 1632.330 906.970 1632.390 ;
        RECT 1084.070 1632.330 1086.970 1632.390 ;
        RECT 1264.070 1632.330 1266.970 1632.390 ;
        RECT 1444.070 1632.330 1446.970 1632.390 ;
        RECT 1624.070 1632.330 1626.970 1632.390 ;
        RECT 1804.070 1632.330 1806.970 1632.390 ;
        RECT 1984.070 1632.330 1986.970 1632.390 ;
        RECT 2164.070 1632.330 2166.970 1632.390 ;
        RECT 2344.070 1632.330 2346.970 1632.390 ;
        RECT 2524.070 1632.330 2526.970 1632.390 ;
        RECT 2704.070 1632.330 2706.970 1632.390 ;
        RECT 2884.070 1632.330 2886.970 1632.390 ;
        RECT 2926.650 1632.330 2929.550 1632.390 ;
        RECT -14.530 1629.430 2934.150 1632.330 ;
        RECT -9.930 1629.370 -7.030 1629.430 ;
        RECT 4.070 1629.370 6.970 1629.430 ;
        RECT 184.070 1629.370 186.970 1629.430 ;
        RECT 364.070 1629.370 366.970 1629.430 ;
        RECT 544.070 1629.370 546.970 1629.430 ;
        RECT 724.070 1629.370 726.970 1629.430 ;
        RECT 904.070 1629.370 906.970 1629.430 ;
        RECT 1084.070 1629.370 1086.970 1629.430 ;
        RECT 1264.070 1629.370 1266.970 1629.430 ;
        RECT 1444.070 1629.370 1446.970 1629.430 ;
        RECT 1624.070 1629.370 1626.970 1629.430 ;
        RECT 1804.070 1629.370 1806.970 1629.430 ;
        RECT 1984.070 1629.370 1986.970 1629.430 ;
        RECT 2164.070 1629.370 2166.970 1629.430 ;
        RECT 2344.070 1629.370 2346.970 1629.430 ;
        RECT 2524.070 1629.370 2526.970 1629.430 ;
        RECT 2704.070 1629.370 2706.970 1629.430 ;
        RECT 2884.070 1629.370 2886.970 1629.430 ;
        RECT 2926.650 1629.370 2929.550 1629.430 ;
        RECT -9.930 1452.330 -7.030 1452.390 ;
        RECT 4.070 1452.330 6.970 1452.390 ;
        RECT 184.070 1452.330 186.970 1452.390 ;
        RECT 364.070 1452.330 366.970 1452.390 ;
        RECT 544.070 1452.330 546.970 1452.390 ;
        RECT 724.070 1452.330 726.970 1452.390 ;
        RECT 904.070 1452.330 906.970 1452.390 ;
        RECT 1084.070 1452.330 1086.970 1452.390 ;
        RECT 1264.070 1452.330 1266.970 1452.390 ;
        RECT 1444.070 1452.330 1446.970 1452.390 ;
        RECT 1624.070 1452.330 1626.970 1452.390 ;
        RECT 1804.070 1452.330 1806.970 1452.390 ;
        RECT 1984.070 1452.330 1986.970 1452.390 ;
        RECT 2164.070 1452.330 2166.970 1452.390 ;
        RECT 2344.070 1452.330 2346.970 1452.390 ;
        RECT 2524.070 1452.330 2526.970 1452.390 ;
        RECT 2704.070 1452.330 2706.970 1452.390 ;
        RECT 2884.070 1452.330 2886.970 1452.390 ;
        RECT 2926.650 1452.330 2929.550 1452.390 ;
        RECT -14.530 1449.430 2934.150 1452.330 ;
        RECT -9.930 1449.370 -7.030 1449.430 ;
        RECT 4.070 1449.370 6.970 1449.430 ;
        RECT 184.070 1449.370 186.970 1449.430 ;
        RECT 364.070 1449.370 366.970 1449.430 ;
        RECT 544.070 1449.370 546.970 1449.430 ;
        RECT 724.070 1449.370 726.970 1449.430 ;
        RECT 904.070 1449.370 906.970 1449.430 ;
        RECT 1084.070 1449.370 1086.970 1449.430 ;
        RECT 1264.070 1449.370 1266.970 1449.430 ;
        RECT 1444.070 1449.370 1446.970 1449.430 ;
        RECT 1624.070 1449.370 1626.970 1449.430 ;
        RECT 1804.070 1449.370 1806.970 1449.430 ;
        RECT 1984.070 1449.370 1986.970 1449.430 ;
        RECT 2164.070 1449.370 2166.970 1449.430 ;
        RECT 2344.070 1449.370 2346.970 1449.430 ;
        RECT 2524.070 1449.370 2526.970 1449.430 ;
        RECT 2704.070 1449.370 2706.970 1449.430 ;
        RECT 2884.070 1449.370 2886.970 1449.430 ;
        RECT 2926.650 1449.370 2929.550 1449.430 ;
        RECT -9.930 1272.330 -7.030 1272.390 ;
        RECT 4.070 1272.330 6.970 1272.390 ;
        RECT 184.070 1272.330 186.970 1272.390 ;
        RECT 364.070 1272.330 366.970 1272.390 ;
        RECT 544.070 1272.330 546.970 1272.390 ;
        RECT 724.070 1272.330 726.970 1272.390 ;
        RECT 904.070 1272.330 906.970 1272.390 ;
        RECT 1084.070 1272.330 1086.970 1272.390 ;
        RECT 1264.070 1272.330 1266.970 1272.390 ;
        RECT 1444.070 1272.330 1446.970 1272.390 ;
        RECT 1624.070 1272.330 1626.970 1272.390 ;
        RECT 1804.070 1272.330 1806.970 1272.390 ;
        RECT 1984.070 1272.330 1986.970 1272.390 ;
        RECT 2164.070 1272.330 2166.970 1272.390 ;
        RECT 2344.070 1272.330 2346.970 1272.390 ;
        RECT 2524.070 1272.330 2526.970 1272.390 ;
        RECT 2704.070 1272.330 2706.970 1272.390 ;
        RECT 2884.070 1272.330 2886.970 1272.390 ;
        RECT 2926.650 1272.330 2929.550 1272.390 ;
        RECT -14.530 1269.430 2934.150 1272.330 ;
        RECT -9.930 1269.370 -7.030 1269.430 ;
        RECT 4.070 1269.370 6.970 1269.430 ;
        RECT 184.070 1269.370 186.970 1269.430 ;
        RECT 364.070 1269.370 366.970 1269.430 ;
        RECT 544.070 1269.370 546.970 1269.430 ;
        RECT 724.070 1269.370 726.970 1269.430 ;
        RECT 904.070 1269.370 906.970 1269.430 ;
        RECT 1084.070 1269.370 1086.970 1269.430 ;
        RECT 1264.070 1269.370 1266.970 1269.430 ;
        RECT 1444.070 1269.370 1446.970 1269.430 ;
        RECT 1624.070 1269.370 1626.970 1269.430 ;
        RECT 1804.070 1269.370 1806.970 1269.430 ;
        RECT 1984.070 1269.370 1986.970 1269.430 ;
        RECT 2164.070 1269.370 2166.970 1269.430 ;
        RECT 2344.070 1269.370 2346.970 1269.430 ;
        RECT 2524.070 1269.370 2526.970 1269.430 ;
        RECT 2704.070 1269.370 2706.970 1269.430 ;
        RECT 2884.070 1269.370 2886.970 1269.430 ;
        RECT 2926.650 1269.370 2929.550 1269.430 ;
        RECT -9.930 1092.330 -7.030 1092.390 ;
        RECT 4.070 1092.330 6.970 1092.390 ;
        RECT 184.070 1092.330 186.970 1092.390 ;
        RECT 364.070 1092.330 366.970 1092.390 ;
        RECT 544.070 1092.330 546.970 1092.390 ;
        RECT 724.070 1092.330 726.970 1092.390 ;
        RECT 904.070 1092.330 906.970 1092.390 ;
        RECT 1084.070 1092.330 1086.970 1092.390 ;
        RECT 1264.070 1092.330 1266.970 1092.390 ;
        RECT 1444.070 1092.330 1446.970 1092.390 ;
        RECT 1624.070 1092.330 1626.970 1092.390 ;
        RECT 1804.070 1092.330 1806.970 1092.390 ;
        RECT 1984.070 1092.330 1986.970 1092.390 ;
        RECT 2164.070 1092.330 2166.970 1092.390 ;
        RECT 2344.070 1092.330 2346.970 1092.390 ;
        RECT 2524.070 1092.330 2526.970 1092.390 ;
        RECT 2704.070 1092.330 2706.970 1092.390 ;
        RECT 2884.070 1092.330 2886.970 1092.390 ;
        RECT 2926.650 1092.330 2929.550 1092.390 ;
        RECT -14.530 1089.430 2934.150 1092.330 ;
        RECT -9.930 1089.370 -7.030 1089.430 ;
        RECT 4.070 1089.370 6.970 1089.430 ;
        RECT 184.070 1089.370 186.970 1089.430 ;
        RECT 364.070 1089.370 366.970 1089.430 ;
        RECT 544.070 1089.370 546.970 1089.430 ;
        RECT 724.070 1089.370 726.970 1089.430 ;
        RECT 904.070 1089.370 906.970 1089.430 ;
        RECT 1084.070 1089.370 1086.970 1089.430 ;
        RECT 1264.070 1089.370 1266.970 1089.430 ;
        RECT 1444.070 1089.370 1446.970 1089.430 ;
        RECT 1624.070 1089.370 1626.970 1089.430 ;
        RECT 1804.070 1089.370 1806.970 1089.430 ;
        RECT 1984.070 1089.370 1986.970 1089.430 ;
        RECT 2164.070 1089.370 2166.970 1089.430 ;
        RECT 2344.070 1089.370 2346.970 1089.430 ;
        RECT 2524.070 1089.370 2526.970 1089.430 ;
        RECT 2704.070 1089.370 2706.970 1089.430 ;
        RECT 2884.070 1089.370 2886.970 1089.430 ;
        RECT 2926.650 1089.370 2929.550 1089.430 ;
        RECT -9.930 912.330 -7.030 912.390 ;
        RECT 4.070 912.330 6.970 912.390 ;
        RECT 184.070 912.330 186.970 912.390 ;
        RECT 364.070 912.330 366.970 912.390 ;
        RECT 544.070 912.330 546.970 912.390 ;
        RECT 724.070 912.330 726.970 912.390 ;
        RECT 904.070 912.330 906.970 912.390 ;
        RECT 1084.070 912.330 1086.970 912.390 ;
        RECT 1264.070 912.330 1266.970 912.390 ;
        RECT 1444.070 912.330 1446.970 912.390 ;
        RECT 1624.070 912.330 1626.970 912.390 ;
        RECT 1804.070 912.330 1806.970 912.390 ;
        RECT 1984.070 912.330 1986.970 912.390 ;
        RECT 2164.070 912.330 2166.970 912.390 ;
        RECT 2344.070 912.330 2346.970 912.390 ;
        RECT 2524.070 912.330 2526.970 912.390 ;
        RECT 2704.070 912.330 2706.970 912.390 ;
        RECT 2884.070 912.330 2886.970 912.390 ;
        RECT 2926.650 912.330 2929.550 912.390 ;
        RECT -14.530 909.430 2934.150 912.330 ;
        RECT -9.930 909.370 -7.030 909.430 ;
        RECT 4.070 909.370 6.970 909.430 ;
        RECT 184.070 909.370 186.970 909.430 ;
        RECT 364.070 909.370 366.970 909.430 ;
        RECT 544.070 909.370 546.970 909.430 ;
        RECT 724.070 909.370 726.970 909.430 ;
        RECT 904.070 909.370 906.970 909.430 ;
        RECT 1084.070 909.370 1086.970 909.430 ;
        RECT 1264.070 909.370 1266.970 909.430 ;
        RECT 1444.070 909.370 1446.970 909.430 ;
        RECT 1624.070 909.370 1626.970 909.430 ;
        RECT 1804.070 909.370 1806.970 909.430 ;
        RECT 1984.070 909.370 1986.970 909.430 ;
        RECT 2164.070 909.370 2166.970 909.430 ;
        RECT 2344.070 909.370 2346.970 909.430 ;
        RECT 2524.070 909.370 2526.970 909.430 ;
        RECT 2704.070 909.370 2706.970 909.430 ;
        RECT 2884.070 909.370 2886.970 909.430 ;
        RECT 2926.650 909.370 2929.550 909.430 ;
        RECT -9.930 732.330 -7.030 732.390 ;
        RECT 4.070 732.330 6.970 732.390 ;
        RECT 184.070 732.330 186.970 732.390 ;
        RECT 364.070 732.330 366.970 732.390 ;
        RECT 544.070 732.330 546.970 732.390 ;
        RECT 724.070 732.330 726.970 732.390 ;
        RECT 904.070 732.330 906.970 732.390 ;
        RECT 1084.070 732.330 1086.970 732.390 ;
        RECT 1264.070 732.330 1266.970 732.390 ;
        RECT 1444.070 732.330 1446.970 732.390 ;
        RECT 1624.070 732.330 1626.970 732.390 ;
        RECT 1804.070 732.330 1806.970 732.390 ;
        RECT 1984.070 732.330 1986.970 732.390 ;
        RECT 2164.070 732.330 2166.970 732.390 ;
        RECT 2344.070 732.330 2346.970 732.390 ;
        RECT 2524.070 732.330 2526.970 732.390 ;
        RECT 2704.070 732.330 2706.970 732.390 ;
        RECT 2884.070 732.330 2886.970 732.390 ;
        RECT 2926.650 732.330 2929.550 732.390 ;
        RECT -14.530 729.430 2934.150 732.330 ;
        RECT -9.930 729.370 -7.030 729.430 ;
        RECT 4.070 729.370 6.970 729.430 ;
        RECT 184.070 729.370 186.970 729.430 ;
        RECT 364.070 729.370 366.970 729.430 ;
        RECT 544.070 729.370 546.970 729.430 ;
        RECT 724.070 729.370 726.970 729.430 ;
        RECT 904.070 729.370 906.970 729.430 ;
        RECT 1084.070 729.370 1086.970 729.430 ;
        RECT 1264.070 729.370 1266.970 729.430 ;
        RECT 1444.070 729.370 1446.970 729.430 ;
        RECT 1624.070 729.370 1626.970 729.430 ;
        RECT 1804.070 729.370 1806.970 729.430 ;
        RECT 1984.070 729.370 1986.970 729.430 ;
        RECT 2164.070 729.370 2166.970 729.430 ;
        RECT 2344.070 729.370 2346.970 729.430 ;
        RECT 2524.070 729.370 2526.970 729.430 ;
        RECT 2704.070 729.370 2706.970 729.430 ;
        RECT 2884.070 729.370 2886.970 729.430 ;
        RECT 2926.650 729.370 2929.550 729.430 ;
        RECT -9.930 552.330 -7.030 552.390 ;
        RECT 4.070 552.330 6.970 552.390 ;
        RECT 184.070 552.330 186.970 552.390 ;
        RECT 364.070 552.330 366.970 552.390 ;
        RECT 544.070 552.330 546.970 552.390 ;
        RECT 724.070 552.330 726.970 552.390 ;
        RECT 904.070 552.330 906.970 552.390 ;
        RECT 1084.070 552.330 1086.970 552.390 ;
        RECT 1264.070 552.330 1266.970 552.390 ;
        RECT 1444.070 552.330 1446.970 552.390 ;
        RECT 1624.070 552.330 1626.970 552.390 ;
        RECT 1804.070 552.330 1806.970 552.390 ;
        RECT 1984.070 552.330 1986.970 552.390 ;
        RECT 2164.070 552.330 2166.970 552.390 ;
        RECT 2344.070 552.330 2346.970 552.390 ;
        RECT 2524.070 552.330 2526.970 552.390 ;
        RECT 2704.070 552.330 2706.970 552.390 ;
        RECT 2884.070 552.330 2886.970 552.390 ;
        RECT 2926.650 552.330 2929.550 552.390 ;
        RECT -14.530 549.430 2934.150 552.330 ;
        RECT -9.930 549.370 -7.030 549.430 ;
        RECT 4.070 549.370 6.970 549.430 ;
        RECT 184.070 549.370 186.970 549.430 ;
        RECT 364.070 549.370 366.970 549.430 ;
        RECT 544.070 549.370 546.970 549.430 ;
        RECT 724.070 549.370 726.970 549.430 ;
        RECT 904.070 549.370 906.970 549.430 ;
        RECT 1084.070 549.370 1086.970 549.430 ;
        RECT 1264.070 549.370 1266.970 549.430 ;
        RECT 1444.070 549.370 1446.970 549.430 ;
        RECT 1624.070 549.370 1626.970 549.430 ;
        RECT 1804.070 549.370 1806.970 549.430 ;
        RECT 1984.070 549.370 1986.970 549.430 ;
        RECT 2164.070 549.370 2166.970 549.430 ;
        RECT 2344.070 549.370 2346.970 549.430 ;
        RECT 2524.070 549.370 2526.970 549.430 ;
        RECT 2704.070 549.370 2706.970 549.430 ;
        RECT 2884.070 549.370 2886.970 549.430 ;
        RECT 2926.650 549.370 2929.550 549.430 ;
        RECT -9.930 372.330 -7.030 372.390 ;
        RECT 4.070 372.330 6.970 372.390 ;
        RECT 184.070 372.330 186.970 372.390 ;
        RECT 364.070 372.330 366.970 372.390 ;
        RECT 544.070 372.330 546.970 372.390 ;
        RECT 724.070 372.330 726.970 372.390 ;
        RECT 904.070 372.330 906.970 372.390 ;
        RECT 1084.070 372.330 1086.970 372.390 ;
        RECT 1264.070 372.330 1266.970 372.390 ;
        RECT 1444.070 372.330 1446.970 372.390 ;
        RECT 1624.070 372.330 1626.970 372.390 ;
        RECT 1804.070 372.330 1806.970 372.390 ;
        RECT 1984.070 372.330 1986.970 372.390 ;
        RECT 2164.070 372.330 2166.970 372.390 ;
        RECT 2344.070 372.330 2346.970 372.390 ;
        RECT 2524.070 372.330 2526.970 372.390 ;
        RECT 2704.070 372.330 2706.970 372.390 ;
        RECT 2884.070 372.330 2886.970 372.390 ;
        RECT 2926.650 372.330 2929.550 372.390 ;
        RECT -14.530 369.430 2934.150 372.330 ;
        RECT -9.930 369.370 -7.030 369.430 ;
        RECT 4.070 369.370 6.970 369.430 ;
        RECT 184.070 369.370 186.970 369.430 ;
        RECT 364.070 369.370 366.970 369.430 ;
        RECT 544.070 369.370 546.970 369.430 ;
        RECT 724.070 369.370 726.970 369.430 ;
        RECT 904.070 369.370 906.970 369.430 ;
        RECT 1084.070 369.370 1086.970 369.430 ;
        RECT 1264.070 369.370 1266.970 369.430 ;
        RECT 1444.070 369.370 1446.970 369.430 ;
        RECT 1624.070 369.370 1626.970 369.430 ;
        RECT 1804.070 369.370 1806.970 369.430 ;
        RECT 1984.070 369.370 1986.970 369.430 ;
        RECT 2164.070 369.370 2166.970 369.430 ;
        RECT 2344.070 369.370 2346.970 369.430 ;
        RECT 2524.070 369.370 2526.970 369.430 ;
        RECT 2704.070 369.370 2706.970 369.430 ;
        RECT 2884.070 369.370 2886.970 369.430 ;
        RECT 2926.650 369.370 2929.550 369.430 ;
        RECT -9.930 192.330 -7.030 192.390 ;
        RECT 4.070 192.330 6.970 192.390 ;
        RECT 184.070 192.330 186.970 192.390 ;
        RECT 364.070 192.330 366.970 192.390 ;
        RECT 544.070 192.330 546.970 192.390 ;
        RECT 724.070 192.330 726.970 192.390 ;
        RECT 904.070 192.330 906.970 192.390 ;
        RECT 1084.070 192.330 1086.970 192.390 ;
        RECT 1264.070 192.330 1266.970 192.390 ;
        RECT 1444.070 192.330 1446.970 192.390 ;
        RECT 1624.070 192.330 1626.970 192.390 ;
        RECT 1804.070 192.330 1806.970 192.390 ;
        RECT 1984.070 192.330 1986.970 192.390 ;
        RECT 2164.070 192.330 2166.970 192.390 ;
        RECT 2344.070 192.330 2346.970 192.390 ;
        RECT 2524.070 192.330 2526.970 192.390 ;
        RECT 2704.070 192.330 2706.970 192.390 ;
        RECT 2884.070 192.330 2886.970 192.390 ;
        RECT 2926.650 192.330 2929.550 192.390 ;
        RECT -14.530 189.430 2934.150 192.330 ;
        RECT -9.930 189.370 -7.030 189.430 ;
        RECT 4.070 189.370 6.970 189.430 ;
        RECT 184.070 189.370 186.970 189.430 ;
        RECT 364.070 189.370 366.970 189.430 ;
        RECT 544.070 189.370 546.970 189.430 ;
        RECT 724.070 189.370 726.970 189.430 ;
        RECT 904.070 189.370 906.970 189.430 ;
        RECT 1084.070 189.370 1086.970 189.430 ;
        RECT 1264.070 189.370 1266.970 189.430 ;
        RECT 1444.070 189.370 1446.970 189.430 ;
        RECT 1624.070 189.370 1626.970 189.430 ;
        RECT 1804.070 189.370 1806.970 189.430 ;
        RECT 1984.070 189.370 1986.970 189.430 ;
        RECT 2164.070 189.370 2166.970 189.430 ;
        RECT 2344.070 189.370 2346.970 189.430 ;
        RECT 2524.070 189.370 2526.970 189.430 ;
        RECT 2704.070 189.370 2706.970 189.430 ;
        RECT 2884.070 189.370 2886.970 189.430 ;
        RECT 2926.650 189.370 2929.550 189.430 ;
        RECT -9.930 12.330 -7.030 12.390 ;
        RECT 4.070 12.330 6.970 12.390 ;
        RECT 184.070 12.330 186.970 12.390 ;
        RECT 364.070 12.330 366.970 12.390 ;
        RECT 544.070 12.330 546.970 12.390 ;
        RECT 724.070 12.330 726.970 12.390 ;
        RECT 904.070 12.330 906.970 12.390 ;
        RECT 1084.070 12.330 1086.970 12.390 ;
        RECT 1264.070 12.330 1266.970 12.390 ;
        RECT 1444.070 12.330 1446.970 12.390 ;
        RECT 1624.070 12.330 1626.970 12.390 ;
        RECT 1804.070 12.330 1806.970 12.390 ;
        RECT 1984.070 12.330 1986.970 12.390 ;
        RECT 2164.070 12.330 2166.970 12.390 ;
        RECT 2344.070 12.330 2346.970 12.390 ;
        RECT 2524.070 12.330 2526.970 12.390 ;
        RECT 2704.070 12.330 2706.970 12.390 ;
        RECT 2884.070 12.330 2886.970 12.390 ;
        RECT 2926.650 12.330 2929.550 12.390 ;
        RECT -14.530 9.430 2934.150 12.330 ;
        RECT -9.930 9.370 -7.030 9.430 ;
        RECT 4.070 9.370 6.970 9.430 ;
        RECT 184.070 9.370 186.970 9.430 ;
        RECT 364.070 9.370 366.970 9.430 ;
        RECT 544.070 9.370 546.970 9.430 ;
        RECT 724.070 9.370 726.970 9.430 ;
        RECT 904.070 9.370 906.970 9.430 ;
        RECT 1084.070 9.370 1086.970 9.430 ;
        RECT 1264.070 9.370 1266.970 9.430 ;
        RECT 1444.070 9.370 1446.970 9.430 ;
        RECT 1624.070 9.370 1626.970 9.430 ;
        RECT 1804.070 9.370 1806.970 9.430 ;
        RECT 1984.070 9.370 1986.970 9.430 ;
        RECT 2164.070 9.370 2166.970 9.430 ;
        RECT 2344.070 9.370 2346.970 9.430 ;
        RECT 2524.070 9.370 2526.970 9.430 ;
        RECT 2704.070 9.370 2706.970 9.430 ;
        RECT 2884.070 9.370 2886.970 9.430 ;
        RECT 2926.650 9.370 2929.550 9.430 ;
        RECT -9.930 -1.670 -7.030 -1.610 ;
        RECT 4.070 -1.670 6.970 -1.610 ;
        RECT 184.070 -1.670 186.970 -1.610 ;
        RECT 364.070 -1.670 366.970 -1.610 ;
        RECT 544.070 -1.670 546.970 -1.610 ;
        RECT 724.070 -1.670 726.970 -1.610 ;
        RECT 904.070 -1.670 906.970 -1.610 ;
        RECT 1084.070 -1.670 1086.970 -1.610 ;
        RECT 1264.070 -1.670 1266.970 -1.610 ;
        RECT 1444.070 -1.670 1446.970 -1.610 ;
        RECT 1624.070 -1.670 1626.970 -1.610 ;
        RECT 1804.070 -1.670 1806.970 -1.610 ;
        RECT 1984.070 -1.670 1986.970 -1.610 ;
        RECT 2164.070 -1.670 2166.970 -1.610 ;
        RECT 2344.070 -1.670 2346.970 -1.610 ;
        RECT 2524.070 -1.670 2526.970 -1.610 ;
        RECT 2704.070 -1.670 2706.970 -1.610 ;
        RECT 2884.070 -1.670 2886.970 -1.610 ;
        RECT 2926.650 -1.670 2929.550 -1.610 ;
        RECT -9.930 -4.570 2929.550 -1.670 ;
        RECT -9.930 -4.630 -7.030 -4.570 ;
        RECT 4.070 -4.630 6.970 -4.570 ;
        RECT 184.070 -4.630 186.970 -4.570 ;
        RECT 364.070 -4.630 366.970 -4.570 ;
        RECT 544.070 -4.630 546.970 -4.570 ;
        RECT 724.070 -4.630 726.970 -4.570 ;
        RECT 904.070 -4.630 906.970 -4.570 ;
        RECT 1084.070 -4.630 1086.970 -4.570 ;
        RECT 1264.070 -4.630 1266.970 -4.570 ;
        RECT 1444.070 -4.630 1446.970 -4.570 ;
        RECT 1624.070 -4.630 1626.970 -4.570 ;
        RECT 1804.070 -4.630 1806.970 -4.570 ;
        RECT 1984.070 -4.630 1986.970 -4.570 ;
        RECT 2164.070 -4.630 2166.970 -4.570 ;
        RECT 2344.070 -4.630 2346.970 -4.570 ;
        RECT 2524.070 -4.630 2526.970 -4.570 ;
        RECT 2704.070 -4.630 2706.970 -4.570 ;
        RECT 2884.070 -4.630 2886.970 -4.570 ;
        RECT 2926.650 -4.630 2929.550 -4.570 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.530 -9.170 -11.630 3528.850 ;
        RECT 94.070 -9.170 96.970 3528.850 ;
        RECT 274.070 -9.170 276.970 3528.850 ;
        RECT 454.070 -9.170 456.970 3528.850 ;
        RECT 634.070 -9.170 636.970 3528.850 ;
        RECT 814.070 -9.170 816.970 3528.850 ;
        RECT 994.070 -9.170 996.970 3528.850 ;
        RECT 1174.070 -9.170 1176.970 3528.850 ;
        RECT 1354.070 -9.170 1356.970 3528.850 ;
        RECT 1534.070 -9.170 1536.970 3528.850 ;
        RECT 1714.070 -9.170 1716.970 3528.850 ;
        RECT 1894.070 -9.170 1896.970 3528.850 ;
        RECT 2074.070 -9.170 2076.970 3528.850 ;
        RECT 2254.070 -9.170 2256.970 3528.850 ;
        RECT 2434.070 -9.170 2436.970 3528.850 ;
        RECT 2614.070 -9.170 2616.970 3528.850 ;
        RECT 2794.070 -9.170 2796.970 3528.850 ;
        RECT 2931.250 -9.170 2934.150 3528.850 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.530 3528.850 -11.630 3528.910 ;
        RECT 94.070 3528.850 96.970 3528.910 ;
        RECT 274.070 3528.850 276.970 3528.910 ;
        RECT 454.070 3528.850 456.970 3528.910 ;
        RECT 634.070 3528.850 636.970 3528.910 ;
        RECT 814.070 3528.850 816.970 3528.910 ;
        RECT 994.070 3528.850 996.970 3528.910 ;
        RECT 1174.070 3528.850 1176.970 3528.910 ;
        RECT 1354.070 3528.850 1356.970 3528.910 ;
        RECT 1534.070 3528.850 1536.970 3528.910 ;
        RECT 1714.070 3528.850 1716.970 3528.910 ;
        RECT 1894.070 3528.850 1896.970 3528.910 ;
        RECT 2074.070 3528.850 2076.970 3528.910 ;
        RECT 2254.070 3528.850 2256.970 3528.910 ;
        RECT 2434.070 3528.850 2436.970 3528.910 ;
        RECT 2614.070 3528.850 2616.970 3528.910 ;
        RECT 2794.070 3528.850 2796.970 3528.910 ;
        RECT 2931.250 3528.850 2934.150 3528.910 ;
        RECT -14.530 3525.950 2934.150 3528.850 ;
        RECT -14.530 3525.890 -11.630 3525.950 ;
        RECT 94.070 3525.890 96.970 3525.950 ;
        RECT 274.070 3525.890 276.970 3525.950 ;
        RECT 454.070 3525.890 456.970 3525.950 ;
        RECT 634.070 3525.890 636.970 3525.950 ;
        RECT 814.070 3525.890 816.970 3525.950 ;
        RECT 994.070 3525.890 996.970 3525.950 ;
        RECT 1174.070 3525.890 1176.970 3525.950 ;
        RECT 1354.070 3525.890 1356.970 3525.950 ;
        RECT 1534.070 3525.890 1536.970 3525.950 ;
        RECT 1714.070 3525.890 1716.970 3525.950 ;
        RECT 1894.070 3525.890 1896.970 3525.950 ;
        RECT 2074.070 3525.890 2076.970 3525.950 ;
        RECT 2254.070 3525.890 2256.970 3525.950 ;
        RECT 2434.070 3525.890 2436.970 3525.950 ;
        RECT 2614.070 3525.890 2616.970 3525.950 ;
        RECT 2794.070 3525.890 2796.970 3525.950 ;
        RECT 2931.250 3525.890 2934.150 3525.950 ;
        RECT -14.530 3342.330 -11.630 3342.390 ;
        RECT 94.070 3342.330 96.970 3342.390 ;
        RECT 274.070 3342.330 276.970 3342.390 ;
        RECT 454.070 3342.330 456.970 3342.390 ;
        RECT 634.070 3342.330 636.970 3342.390 ;
        RECT 814.070 3342.330 816.970 3342.390 ;
        RECT 994.070 3342.330 996.970 3342.390 ;
        RECT 1174.070 3342.330 1176.970 3342.390 ;
        RECT 1354.070 3342.330 1356.970 3342.390 ;
        RECT 1534.070 3342.330 1536.970 3342.390 ;
        RECT 1714.070 3342.330 1716.970 3342.390 ;
        RECT 1894.070 3342.330 1896.970 3342.390 ;
        RECT 2074.070 3342.330 2076.970 3342.390 ;
        RECT 2254.070 3342.330 2256.970 3342.390 ;
        RECT 2434.070 3342.330 2436.970 3342.390 ;
        RECT 2614.070 3342.330 2616.970 3342.390 ;
        RECT 2794.070 3342.330 2796.970 3342.390 ;
        RECT 2931.250 3342.330 2934.150 3342.390 ;
        RECT -14.530 3339.430 2934.150 3342.330 ;
        RECT -14.530 3339.370 -11.630 3339.430 ;
        RECT 94.070 3339.370 96.970 3339.430 ;
        RECT 274.070 3339.370 276.970 3339.430 ;
        RECT 454.070 3339.370 456.970 3339.430 ;
        RECT 634.070 3339.370 636.970 3339.430 ;
        RECT 814.070 3339.370 816.970 3339.430 ;
        RECT 994.070 3339.370 996.970 3339.430 ;
        RECT 1174.070 3339.370 1176.970 3339.430 ;
        RECT 1354.070 3339.370 1356.970 3339.430 ;
        RECT 1534.070 3339.370 1536.970 3339.430 ;
        RECT 1714.070 3339.370 1716.970 3339.430 ;
        RECT 1894.070 3339.370 1896.970 3339.430 ;
        RECT 2074.070 3339.370 2076.970 3339.430 ;
        RECT 2254.070 3339.370 2256.970 3339.430 ;
        RECT 2434.070 3339.370 2436.970 3339.430 ;
        RECT 2614.070 3339.370 2616.970 3339.430 ;
        RECT 2794.070 3339.370 2796.970 3339.430 ;
        RECT 2931.250 3339.370 2934.150 3339.430 ;
        RECT -14.530 3162.330 -11.630 3162.390 ;
        RECT 94.070 3162.330 96.970 3162.390 ;
        RECT 274.070 3162.330 276.970 3162.390 ;
        RECT 454.070 3162.330 456.970 3162.390 ;
        RECT 634.070 3162.330 636.970 3162.390 ;
        RECT 814.070 3162.330 816.970 3162.390 ;
        RECT 994.070 3162.330 996.970 3162.390 ;
        RECT 1174.070 3162.330 1176.970 3162.390 ;
        RECT 1354.070 3162.330 1356.970 3162.390 ;
        RECT 1534.070 3162.330 1536.970 3162.390 ;
        RECT 1714.070 3162.330 1716.970 3162.390 ;
        RECT 1894.070 3162.330 1896.970 3162.390 ;
        RECT 2074.070 3162.330 2076.970 3162.390 ;
        RECT 2254.070 3162.330 2256.970 3162.390 ;
        RECT 2434.070 3162.330 2436.970 3162.390 ;
        RECT 2614.070 3162.330 2616.970 3162.390 ;
        RECT 2794.070 3162.330 2796.970 3162.390 ;
        RECT 2931.250 3162.330 2934.150 3162.390 ;
        RECT -14.530 3159.430 2934.150 3162.330 ;
        RECT -14.530 3159.370 -11.630 3159.430 ;
        RECT 94.070 3159.370 96.970 3159.430 ;
        RECT 274.070 3159.370 276.970 3159.430 ;
        RECT 454.070 3159.370 456.970 3159.430 ;
        RECT 634.070 3159.370 636.970 3159.430 ;
        RECT 814.070 3159.370 816.970 3159.430 ;
        RECT 994.070 3159.370 996.970 3159.430 ;
        RECT 1174.070 3159.370 1176.970 3159.430 ;
        RECT 1354.070 3159.370 1356.970 3159.430 ;
        RECT 1534.070 3159.370 1536.970 3159.430 ;
        RECT 1714.070 3159.370 1716.970 3159.430 ;
        RECT 1894.070 3159.370 1896.970 3159.430 ;
        RECT 2074.070 3159.370 2076.970 3159.430 ;
        RECT 2254.070 3159.370 2256.970 3159.430 ;
        RECT 2434.070 3159.370 2436.970 3159.430 ;
        RECT 2614.070 3159.370 2616.970 3159.430 ;
        RECT 2794.070 3159.370 2796.970 3159.430 ;
        RECT 2931.250 3159.370 2934.150 3159.430 ;
        RECT -14.530 2982.330 -11.630 2982.390 ;
        RECT 94.070 2982.330 96.970 2982.390 ;
        RECT 274.070 2982.330 276.970 2982.390 ;
        RECT 454.070 2982.330 456.970 2982.390 ;
        RECT 634.070 2982.330 636.970 2982.390 ;
        RECT 814.070 2982.330 816.970 2982.390 ;
        RECT 994.070 2982.330 996.970 2982.390 ;
        RECT 1174.070 2982.330 1176.970 2982.390 ;
        RECT 1354.070 2982.330 1356.970 2982.390 ;
        RECT 1534.070 2982.330 1536.970 2982.390 ;
        RECT 1714.070 2982.330 1716.970 2982.390 ;
        RECT 1894.070 2982.330 1896.970 2982.390 ;
        RECT 2074.070 2982.330 2076.970 2982.390 ;
        RECT 2254.070 2982.330 2256.970 2982.390 ;
        RECT 2434.070 2982.330 2436.970 2982.390 ;
        RECT 2614.070 2982.330 2616.970 2982.390 ;
        RECT 2794.070 2982.330 2796.970 2982.390 ;
        RECT 2931.250 2982.330 2934.150 2982.390 ;
        RECT -14.530 2979.430 2934.150 2982.330 ;
        RECT -14.530 2979.370 -11.630 2979.430 ;
        RECT 94.070 2979.370 96.970 2979.430 ;
        RECT 274.070 2979.370 276.970 2979.430 ;
        RECT 454.070 2979.370 456.970 2979.430 ;
        RECT 634.070 2979.370 636.970 2979.430 ;
        RECT 814.070 2979.370 816.970 2979.430 ;
        RECT 994.070 2979.370 996.970 2979.430 ;
        RECT 1174.070 2979.370 1176.970 2979.430 ;
        RECT 1354.070 2979.370 1356.970 2979.430 ;
        RECT 1534.070 2979.370 1536.970 2979.430 ;
        RECT 1714.070 2979.370 1716.970 2979.430 ;
        RECT 1894.070 2979.370 1896.970 2979.430 ;
        RECT 2074.070 2979.370 2076.970 2979.430 ;
        RECT 2254.070 2979.370 2256.970 2979.430 ;
        RECT 2434.070 2979.370 2436.970 2979.430 ;
        RECT 2614.070 2979.370 2616.970 2979.430 ;
        RECT 2794.070 2979.370 2796.970 2979.430 ;
        RECT 2931.250 2979.370 2934.150 2979.430 ;
        RECT -14.530 2802.330 -11.630 2802.390 ;
        RECT 94.070 2802.330 96.970 2802.390 ;
        RECT 274.070 2802.330 276.970 2802.390 ;
        RECT 454.070 2802.330 456.970 2802.390 ;
        RECT 634.070 2802.330 636.970 2802.390 ;
        RECT 814.070 2802.330 816.970 2802.390 ;
        RECT 994.070 2802.330 996.970 2802.390 ;
        RECT 1174.070 2802.330 1176.970 2802.390 ;
        RECT 1354.070 2802.330 1356.970 2802.390 ;
        RECT 1534.070 2802.330 1536.970 2802.390 ;
        RECT 1714.070 2802.330 1716.970 2802.390 ;
        RECT 1894.070 2802.330 1896.970 2802.390 ;
        RECT 2074.070 2802.330 2076.970 2802.390 ;
        RECT 2254.070 2802.330 2256.970 2802.390 ;
        RECT 2434.070 2802.330 2436.970 2802.390 ;
        RECT 2614.070 2802.330 2616.970 2802.390 ;
        RECT 2794.070 2802.330 2796.970 2802.390 ;
        RECT 2931.250 2802.330 2934.150 2802.390 ;
        RECT -14.530 2799.430 2934.150 2802.330 ;
        RECT -14.530 2799.370 -11.630 2799.430 ;
        RECT 94.070 2799.370 96.970 2799.430 ;
        RECT 274.070 2799.370 276.970 2799.430 ;
        RECT 454.070 2799.370 456.970 2799.430 ;
        RECT 634.070 2799.370 636.970 2799.430 ;
        RECT 814.070 2799.370 816.970 2799.430 ;
        RECT 994.070 2799.370 996.970 2799.430 ;
        RECT 1174.070 2799.370 1176.970 2799.430 ;
        RECT 1354.070 2799.370 1356.970 2799.430 ;
        RECT 1534.070 2799.370 1536.970 2799.430 ;
        RECT 1714.070 2799.370 1716.970 2799.430 ;
        RECT 1894.070 2799.370 1896.970 2799.430 ;
        RECT 2074.070 2799.370 2076.970 2799.430 ;
        RECT 2254.070 2799.370 2256.970 2799.430 ;
        RECT 2434.070 2799.370 2436.970 2799.430 ;
        RECT 2614.070 2799.370 2616.970 2799.430 ;
        RECT 2794.070 2799.370 2796.970 2799.430 ;
        RECT 2931.250 2799.370 2934.150 2799.430 ;
        RECT -14.530 2622.330 -11.630 2622.390 ;
        RECT 94.070 2622.330 96.970 2622.390 ;
        RECT 274.070 2622.330 276.970 2622.390 ;
        RECT 454.070 2622.330 456.970 2622.390 ;
        RECT 634.070 2622.330 636.970 2622.390 ;
        RECT 814.070 2622.330 816.970 2622.390 ;
        RECT 994.070 2622.330 996.970 2622.390 ;
        RECT 1174.070 2622.330 1176.970 2622.390 ;
        RECT 1354.070 2622.330 1356.970 2622.390 ;
        RECT 1534.070 2622.330 1536.970 2622.390 ;
        RECT 1714.070 2622.330 1716.970 2622.390 ;
        RECT 1894.070 2622.330 1896.970 2622.390 ;
        RECT 2074.070 2622.330 2076.970 2622.390 ;
        RECT 2254.070 2622.330 2256.970 2622.390 ;
        RECT 2434.070 2622.330 2436.970 2622.390 ;
        RECT 2614.070 2622.330 2616.970 2622.390 ;
        RECT 2794.070 2622.330 2796.970 2622.390 ;
        RECT 2931.250 2622.330 2934.150 2622.390 ;
        RECT -14.530 2619.430 2934.150 2622.330 ;
        RECT -14.530 2619.370 -11.630 2619.430 ;
        RECT 94.070 2619.370 96.970 2619.430 ;
        RECT 274.070 2619.370 276.970 2619.430 ;
        RECT 454.070 2619.370 456.970 2619.430 ;
        RECT 634.070 2619.370 636.970 2619.430 ;
        RECT 814.070 2619.370 816.970 2619.430 ;
        RECT 994.070 2619.370 996.970 2619.430 ;
        RECT 1174.070 2619.370 1176.970 2619.430 ;
        RECT 1354.070 2619.370 1356.970 2619.430 ;
        RECT 1534.070 2619.370 1536.970 2619.430 ;
        RECT 1714.070 2619.370 1716.970 2619.430 ;
        RECT 1894.070 2619.370 1896.970 2619.430 ;
        RECT 2074.070 2619.370 2076.970 2619.430 ;
        RECT 2254.070 2619.370 2256.970 2619.430 ;
        RECT 2434.070 2619.370 2436.970 2619.430 ;
        RECT 2614.070 2619.370 2616.970 2619.430 ;
        RECT 2794.070 2619.370 2796.970 2619.430 ;
        RECT 2931.250 2619.370 2934.150 2619.430 ;
        RECT -14.530 2442.330 -11.630 2442.390 ;
        RECT 94.070 2442.330 96.970 2442.390 ;
        RECT 274.070 2442.330 276.970 2442.390 ;
        RECT 454.070 2442.330 456.970 2442.390 ;
        RECT 634.070 2442.330 636.970 2442.390 ;
        RECT 814.070 2442.330 816.970 2442.390 ;
        RECT 994.070 2442.330 996.970 2442.390 ;
        RECT 1174.070 2442.330 1176.970 2442.390 ;
        RECT 1354.070 2442.330 1356.970 2442.390 ;
        RECT 1534.070 2442.330 1536.970 2442.390 ;
        RECT 1714.070 2442.330 1716.970 2442.390 ;
        RECT 1894.070 2442.330 1896.970 2442.390 ;
        RECT 2074.070 2442.330 2076.970 2442.390 ;
        RECT 2254.070 2442.330 2256.970 2442.390 ;
        RECT 2434.070 2442.330 2436.970 2442.390 ;
        RECT 2614.070 2442.330 2616.970 2442.390 ;
        RECT 2794.070 2442.330 2796.970 2442.390 ;
        RECT 2931.250 2442.330 2934.150 2442.390 ;
        RECT -14.530 2439.430 2934.150 2442.330 ;
        RECT -14.530 2439.370 -11.630 2439.430 ;
        RECT 94.070 2439.370 96.970 2439.430 ;
        RECT 274.070 2439.370 276.970 2439.430 ;
        RECT 454.070 2439.370 456.970 2439.430 ;
        RECT 634.070 2439.370 636.970 2439.430 ;
        RECT 814.070 2439.370 816.970 2439.430 ;
        RECT 994.070 2439.370 996.970 2439.430 ;
        RECT 1174.070 2439.370 1176.970 2439.430 ;
        RECT 1354.070 2439.370 1356.970 2439.430 ;
        RECT 1534.070 2439.370 1536.970 2439.430 ;
        RECT 1714.070 2439.370 1716.970 2439.430 ;
        RECT 1894.070 2439.370 1896.970 2439.430 ;
        RECT 2074.070 2439.370 2076.970 2439.430 ;
        RECT 2254.070 2439.370 2256.970 2439.430 ;
        RECT 2434.070 2439.370 2436.970 2439.430 ;
        RECT 2614.070 2439.370 2616.970 2439.430 ;
        RECT 2794.070 2439.370 2796.970 2439.430 ;
        RECT 2931.250 2439.370 2934.150 2439.430 ;
        RECT -14.530 2262.330 -11.630 2262.390 ;
        RECT 94.070 2262.330 96.970 2262.390 ;
        RECT 274.070 2262.330 276.970 2262.390 ;
        RECT 454.070 2262.330 456.970 2262.390 ;
        RECT 634.070 2262.330 636.970 2262.390 ;
        RECT 814.070 2262.330 816.970 2262.390 ;
        RECT 994.070 2262.330 996.970 2262.390 ;
        RECT 1174.070 2262.330 1176.970 2262.390 ;
        RECT 1354.070 2262.330 1356.970 2262.390 ;
        RECT 1534.070 2262.330 1536.970 2262.390 ;
        RECT 1714.070 2262.330 1716.970 2262.390 ;
        RECT 1894.070 2262.330 1896.970 2262.390 ;
        RECT 2074.070 2262.330 2076.970 2262.390 ;
        RECT 2254.070 2262.330 2256.970 2262.390 ;
        RECT 2434.070 2262.330 2436.970 2262.390 ;
        RECT 2614.070 2262.330 2616.970 2262.390 ;
        RECT 2794.070 2262.330 2796.970 2262.390 ;
        RECT 2931.250 2262.330 2934.150 2262.390 ;
        RECT -14.530 2259.430 2934.150 2262.330 ;
        RECT -14.530 2259.370 -11.630 2259.430 ;
        RECT 94.070 2259.370 96.970 2259.430 ;
        RECT 274.070 2259.370 276.970 2259.430 ;
        RECT 454.070 2259.370 456.970 2259.430 ;
        RECT 634.070 2259.370 636.970 2259.430 ;
        RECT 814.070 2259.370 816.970 2259.430 ;
        RECT 994.070 2259.370 996.970 2259.430 ;
        RECT 1174.070 2259.370 1176.970 2259.430 ;
        RECT 1354.070 2259.370 1356.970 2259.430 ;
        RECT 1534.070 2259.370 1536.970 2259.430 ;
        RECT 1714.070 2259.370 1716.970 2259.430 ;
        RECT 1894.070 2259.370 1896.970 2259.430 ;
        RECT 2074.070 2259.370 2076.970 2259.430 ;
        RECT 2254.070 2259.370 2256.970 2259.430 ;
        RECT 2434.070 2259.370 2436.970 2259.430 ;
        RECT 2614.070 2259.370 2616.970 2259.430 ;
        RECT 2794.070 2259.370 2796.970 2259.430 ;
        RECT 2931.250 2259.370 2934.150 2259.430 ;
        RECT -14.530 2082.330 -11.630 2082.390 ;
        RECT 94.070 2082.330 96.970 2082.390 ;
        RECT 274.070 2082.330 276.970 2082.390 ;
        RECT 454.070 2082.330 456.970 2082.390 ;
        RECT 634.070 2082.330 636.970 2082.390 ;
        RECT 814.070 2082.330 816.970 2082.390 ;
        RECT 994.070 2082.330 996.970 2082.390 ;
        RECT 1174.070 2082.330 1176.970 2082.390 ;
        RECT 1354.070 2082.330 1356.970 2082.390 ;
        RECT 1534.070 2082.330 1536.970 2082.390 ;
        RECT 1714.070 2082.330 1716.970 2082.390 ;
        RECT 1894.070 2082.330 1896.970 2082.390 ;
        RECT 2074.070 2082.330 2076.970 2082.390 ;
        RECT 2254.070 2082.330 2256.970 2082.390 ;
        RECT 2434.070 2082.330 2436.970 2082.390 ;
        RECT 2614.070 2082.330 2616.970 2082.390 ;
        RECT 2794.070 2082.330 2796.970 2082.390 ;
        RECT 2931.250 2082.330 2934.150 2082.390 ;
        RECT -14.530 2079.430 2934.150 2082.330 ;
        RECT -14.530 2079.370 -11.630 2079.430 ;
        RECT 94.070 2079.370 96.970 2079.430 ;
        RECT 274.070 2079.370 276.970 2079.430 ;
        RECT 454.070 2079.370 456.970 2079.430 ;
        RECT 634.070 2079.370 636.970 2079.430 ;
        RECT 814.070 2079.370 816.970 2079.430 ;
        RECT 994.070 2079.370 996.970 2079.430 ;
        RECT 1174.070 2079.370 1176.970 2079.430 ;
        RECT 1354.070 2079.370 1356.970 2079.430 ;
        RECT 1534.070 2079.370 1536.970 2079.430 ;
        RECT 1714.070 2079.370 1716.970 2079.430 ;
        RECT 1894.070 2079.370 1896.970 2079.430 ;
        RECT 2074.070 2079.370 2076.970 2079.430 ;
        RECT 2254.070 2079.370 2256.970 2079.430 ;
        RECT 2434.070 2079.370 2436.970 2079.430 ;
        RECT 2614.070 2079.370 2616.970 2079.430 ;
        RECT 2794.070 2079.370 2796.970 2079.430 ;
        RECT 2931.250 2079.370 2934.150 2079.430 ;
        RECT -14.530 1902.330 -11.630 1902.390 ;
        RECT 94.070 1902.330 96.970 1902.390 ;
        RECT 274.070 1902.330 276.970 1902.390 ;
        RECT 454.070 1902.330 456.970 1902.390 ;
        RECT 634.070 1902.330 636.970 1902.390 ;
        RECT 814.070 1902.330 816.970 1902.390 ;
        RECT 994.070 1902.330 996.970 1902.390 ;
        RECT 1174.070 1902.330 1176.970 1902.390 ;
        RECT 1354.070 1902.330 1356.970 1902.390 ;
        RECT 1534.070 1902.330 1536.970 1902.390 ;
        RECT 1714.070 1902.330 1716.970 1902.390 ;
        RECT 1894.070 1902.330 1896.970 1902.390 ;
        RECT 2074.070 1902.330 2076.970 1902.390 ;
        RECT 2254.070 1902.330 2256.970 1902.390 ;
        RECT 2434.070 1902.330 2436.970 1902.390 ;
        RECT 2614.070 1902.330 2616.970 1902.390 ;
        RECT 2794.070 1902.330 2796.970 1902.390 ;
        RECT 2931.250 1902.330 2934.150 1902.390 ;
        RECT -14.530 1899.430 2934.150 1902.330 ;
        RECT -14.530 1899.370 -11.630 1899.430 ;
        RECT 94.070 1899.370 96.970 1899.430 ;
        RECT 274.070 1899.370 276.970 1899.430 ;
        RECT 454.070 1899.370 456.970 1899.430 ;
        RECT 634.070 1899.370 636.970 1899.430 ;
        RECT 814.070 1899.370 816.970 1899.430 ;
        RECT 994.070 1899.370 996.970 1899.430 ;
        RECT 1174.070 1899.370 1176.970 1899.430 ;
        RECT 1354.070 1899.370 1356.970 1899.430 ;
        RECT 1534.070 1899.370 1536.970 1899.430 ;
        RECT 1714.070 1899.370 1716.970 1899.430 ;
        RECT 1894.070 1899.370 1896.970 1899.430 ;
        RECT 2074.070 1899.370 2076.970 1899.430 ;
        RECT 2254.070 1899.370 2256.970 1899.430 ;
        RECT 2434.070 1899.370 2436.970 1899.430 ;
        RECT 2614.070 1899.370 2616.970 1899.430 ;
        RECT 2794.070 1899.370 2796.970 1899.430 ;
        RECT 2931.250 1899.370 2934.150 1899.430 ;
        RECT -14.530 1722.330 -11.630 1722.390 ;
        RECT 94.070 1722.330 96.970 1722.390 ;
        RECT 274.070 1722.330 276.970 1722.390 ;
        RECT 454.070 1722.330 456.970 1722.390 ;
        RECT 634.070 1722.330 636.970 1722.390 ;
        RECT 814.070 1722.330 816.970 1722.390 ;
        RECT 994.070 1722.330 996.970 1722.390 ;
        RECT 1174.070 1722.330 1176.970 1722.390 ;
        RECT 1354.070 1722.330 1356.970 1722.390 ;
        RECT 1534.070 1722.330 1536.970 1722.390 ;
        RECT 1714.070 1722.330 1716.970 1722.390 ;
        RECT 1894.070 1722.330 1896.970 1722.390 ;
        RECT 2074.070 1722.330 2076.970 1722.390 ;
        RECT 2254.070 1722.330 2256.970 1722.390 ;
        RECT 2434.070 1722.330 2436.970 1722.390 ;
        RECT 2614.070 1722.330 2616.970 1722.390 ;
        RECT 2794.070 1722.330 2796.970 1722.390 ;
        RECT 2931.250 1722.330 2934.150 1722.390 ;
        RECT -14.530 1719.430 2934.150 1722.330 ;
        RECT -14.530 1719.370 -11.630 1719.430 ;
        RECT 94.070 1719.370 96.970 1719.430 ;
        RECT 274.070 1719.370 276.970 1719.430 ;
        RECT 454.070 1719.370 456.970 1719.430 ;
        RECT 634.070 1719.370 636.970 1719.430 ;
        RECT 814.070 1719.370 816.970 1719.430 ;
        RECT 994.070 1719.370 996.970 1719.430 ;
        RECT 1174.070 1719.370 1176.970 1719.430 ;
        RECT 1354.070 1719.370 1356.970 1719.430 ;
        RECT 1534.070 1719.370 1536.970 1719.430 ;
        RECT 1714.070 1719.370 1716.970 1719.430 ;
        RECT 1894.070 1719.370 1896.970 1719.430 ;
        RECT 2074.070 1719.370 2076.970 1719.430 ;
        RECT 2254.070 1719.370 2256.970 1719.430 ;
        RECT 2434.070 1719.370 2436.970 1719.430 ;
        RECT 2614.070 1719.370 2616.970 1719.430 ;
        RECT 2794.070 1719.370 2796.970 1719.430 ;
        RECT 2931.250 1719.370 2934.150 1719.430 ;
        RECT -14.530 1542.330 -11.630 1542.390 ;
        RECT 94.070 1542.330 96.970 1542.390 ;
        RECT 274.070 1542.330 276.970 1542.390 ;
        RECT 454.070 1542.330 456.970 1542.390 ;
        RECT 634.070 1542.330 636.970 1542.390 ;
        RECT 814.070 1542.330 816.970 1542.390 ;
        RECT 994.070 1542.330 996.970 1542.390 ;
        RECT 1174.070 1542.330 1176.970 1542.390 ;
        RECT 1354.070 1542.330 1356.970 1542.390 ;
        RECT 1534.070 1542.330 1536.970 1542.390 ;
        RECT 1714.070 1542.330 1716.970 1542.390 ;
        RECT 1894.070 1542.330 1896.970 1542.390 ;
        RECT 2074.070 1542.330 2076.970 1542.390 ;
        RECT 2254.070 1542.330 2256.970 1542.390 ;
        RECT 2434.070 1542.330 2436.970 1542.390 ;
        RECT 2614.070 1542.330 2616.970 1542.390 ;
        RECT 2794.070 1542.330 2796.970 1542.390 ;
        RECT 2931.250 1542.330 2934.150 1542.390 ;
        RECT -14.530 1539.430 2934.150 1542.330 ;
        RECT -14.530 1539.370 -11.630 1539.430 ;
        RECT 94.070 1539.370 96.970 1539.430 ;
        RECT 274.070 1539.370 276.970 1539.430 ;
        RECT 454.070 1539.370 456.970 1539.430 ;
        RECT 634.070 1539.370 636.970 1539.430 ;
        RECT 814.070 1539.370 816.970 1539.430 ;
        RECT 994.070 1539.370 996.970 1539.430 ;
        RECT 1174.070 1539.370 1176.970 1539.430 ;
        RECT 1354.070 1539.370 1356.970 1539.430 ;
        RECT 1534.070 1539.370 1536.970 1539.430 ;
        RECT 1714.070 1539.370 1716.970 1539.430 ;
        RECT 1894.070 1539.370 1896.970 1539.430 ;
        RECT 2074.070 1539.370 2076.970 1539.430 ;
        RECT 2254.070 1539.370 2256.970 1539.430 ;
        RECT 2434.070 1539.370 2436.970 1539.430 ;
        RECT 2614.070 1539.370 2616.970 1539.430 ;
        RECT 2794.070 1539.370 2796.970 1539.430 ;
        RECT 2931.250 1539.370 2934.150 1539.430 ;
        RECT -14.530 1362.330 -11.630 1362.390 ;
        RECT 94.070 1362.330 96.970 1362.390 ;
        RECT 274.070 1362.330 276.970 1362.390 ;
        RECT 454.070 1362.330 456.970 1362.390 ;
        RECT 634.070 1362.330 636.970 1362.390 ;
        RECT 814.070 1362.330 816.970 1362.390 ;
        RECT 994.070 1362.330 996.970 1362.390 ;
        RECT 1174.070 1362.330 1176.970 1362.390 ;
        RECT 1354.070 1362.330 1356.970 1362.390 ;
        RECT 1534.070 1362.330 1536.970 1362.390 ;
        RECT 1714.070 1362.330 1716.970 1362.390 ;
        RECT 1894.070 1362.330 1896.970 1362.390 ;
        RECT 2074.070 1362.330 2076.970 1362.390 ;
        RECT 2254.070 1362.330 2256.970 1362.390 ;
        RECT 2434.070 1362.330 2436.970 1362.390 ;
        RECT 2614.070 1362.330 2616.970 1362.390 ;
        RECT 2794.070 1362.330 2796.970 1362.390 ;
        RECT 2931.250 1362.330 2934.150 1362.390 ;
        RECT -14.530 1359.430 2934.150 1362.330 ;
        RECT -14.530 1359.370 -11.630 1359.430 ;
        RECT 94.070 1359.370 96.970 1359.430 ;
        RECT 274.070 1359.370 276.970 1359.430 ;
        RECT 454.070 1359.370 456.970 1359.430 ;
        RECT 634.070 1359.370 636.970 1359.430 ;
        RECT 814.070 1359.370 816.970 1359.430 ;
        RECT 994.070 1359.370 996.970 1359.430 ;
        RECT 1174.070 1359.370 1176.970 1359.430 ;
        RECT 1354.070 1359.370 1356.970 1359.430 ;
        RECT 1534.070 1359.370 1536.970 1359.430 ;
        RECT 1714.070 1359.370 1716.970 1359.430 ;
        RECT 1894.070 1359.370 1896.970 1359.430 ;
        RECT 2074.070 1359.370 2076.970 1359.430 ;
        RECT 2254.070 1359.370 2256.970 1359.430 ;
        RECT 2434.070 1359.370 2436.970 1359.430 ;
        RECT 2614.070 1359.370 2616.970 1359.430 ;
        RECT 2794.070 1359.370 2796.970 1359.430 ;
        RECT 2931.250 1359.370 2934.150 1359.430 ;
        RECT -14.530 1182.330 -11.630 1182.390 ;
        RECT 94.070 1182.330 96.970 1182.390 ;
        RECT 274.070 1182.330 276.970 1182.390 ;
        RECT 454.070 1182.330 456.970 1182.390 ;
        RECT 634.070 1182.330 636.970 1182.390 ;
        RECT 814.070 1182.330 816.970 1182.390 ;
        RECT 994.070 1182.330 996.970 1182.390 ;
        RECT 1174.070 1182.330 1176.970 1182.390 ;
        RECT 1354.070 1182.330 1356.970 1182.390 ;
        RECT 1534.070 1182.330 1536.970 1182.390 ;
        RECT 1714.070 1182.330 1716.970 1182.390 ;
        RECT 1894.070 1182.330 1896.970 1182.390 ;
        RECT 2074.070 1182.330 2076.970 1182.390 ;
        RECT 2254.070 1182.330 2256.970 1182.390 ;
        RECT 2434.070 1182.330 2436.970 1182.390 ;
        RECT 2614.070 1182.330 2616.970 1182.390 ;
        RECT 2794.070 1182.330 2796.970 1182.390 ;
        RECT 2931.250 1182.330 2934.150 1182.390 ;
        RECT -14.530 1179.430 2934.150 1182.330 ;
        RECT -14.530 1179.370 -11.630 1179.430 ;
        RECT 94.070 1179.370 96.970 1179.430 ;
        RECT 274.070 1179.370 276.970 1179.430 ;
        RECT 454.070 1179.370 456.970 1179.430 ;
        RECT 634.070 1179.370 636.970 1179.430 ;
        RECT 814.070 1179.370 816.970 1179.430 ;
        RECT 994.070 1179.370 996.970 1179.430 ;
        RECT 1174.070 1179.370 1176.970 1179.430 ;
        RECT 1354.070 1179.370 1356.970 1179.430 ;
        RECT 1534.070 1179.370 1536.970 1179.430 ;
        RECT 1714.070 1179.370 1716.970 1179.430 ;
        RECT 1894.070 1179.370 1896.970 1179.430 ;
        RECT 2074.070 1179.370 2076.970 1179.430 ;
        RECT 2254.070 1179.370 2256.970 1179.430 ;
        RECT 2434.070 1179.370 2436.970 1179.430 ;
        RECT 2614.070 1179.370 2616.970 1179.430 ;
        RECT 2794.070 1179.370 2796.970 1179.430 ;
        RECT 2931.250 1179.370 2934.150 1179.430 ;
        RECT -14.530 1002.330 -11.630 1002.390 ;
        RECT 94.070 1002.330 96.970 1002.390 ;
        RECT 274.070 1002.330 276.970 1002.390 ;
        RECT 454.070 1002.330 456.970 1002.390 ;
        RECT 634.070 1002.330 636.970 1002.390 ;
        RECT 814.070 1002.330 816.970 1002.390 ;
        RECT 994.070 1002.330 996.970 1002.390 ;
        RECT 1174.070 1002.330 1176.970 1002.390 ;
        RECT 1354.070 1002.330 1356.970 1002.390 ;
        RECT 1534.070 1002.330 1536.970 1002.390 ;
        RECT 1714.070 1002.330 1716.970 1002.390 ;
        RECT 1894.070 1002.330 1896.970 1002.390 ;
        RECT 2074.070 1002.330 2076.970 1002.390 ;
        RECT 2254.070 1002.330 2256.970 1002.390 ;
        RECT 2434.070 1002.330 2436.970 1002.390 ;
        RECT 2614.070 1002.330 2616.970 1002.390 ;
        RECT 2794.070 1002.330 2796.970 1002.390 ;
        RECT 2931.250 1002.330 2934.150 1002.390 ;
        RECT -14.530 999.430 2934.150 1002.330 ;
        RECT -14.530 999.370 -11.630 999.430 ;
        RECT 94.070 999.370 96.970 999.430 ;
        RECT 274.070 999.370 276.970 999.430 ;
        RECT 454.070 999.370 456.970 999.430 ;
        RECT 634.070 999.370 636.970 999.430 ;
        RECT 814.070 999.370 816.970 999.430 ;
        RECT 994.070 999.370 996.970 999.430 ;
        RECT 1174.070 999.370 1176.970 999.430 ;
        RECT 1354.070 999.370 1356.970 999.430 ;
        RECT 1534.070 999.370 1536.970 999.430 ;
        RECT 1714.070 999.370 1716.970 999.430 ;
        RECT 1894.070 999.370 1896.970 999.430 ;
        RECT 2074.070 999.370 2076.970 999.430 ;
        RECT 2254.070 999.370 2256.970 999.430 ;
        RECT 2434.070 999.370 2436.970 999.430 ;
        RECT 2614.070 999.370 2616.970 999.430 ;
        RECT 2794.070 999.370 2796.970 999.430 ;
        RECT 2931.250 999.370 2934.150 999.430 ;
        RECT -14.530 822.330 -11.630 822.390 ;
        RECT 94.070 822.330 96.970 822.390 ;
        RECT 274.070 822.330 276.970 822.390 ;
        RECT 454.070 822.330 456.970 822.390 ;
        RECT 634.070 822.330 636.970 822.390 ;
        RECT 814.070 822.330 816.970 822.390 ;
        RECT 994.070 822.330 996.970 822.390 ;
        RECT 1174.070 822.330 1176.970 822.390 ;
        RECT 1354.070 822.330 1356.970 822.390 ;
        RECT 1534.070 822.330 1536.970 822.390 ;
        RECT 1714.070 822.330 1716.970 822.390 ;
        RECT 1894.070 822.330 1896.970 822.390 ;
        RECT 2074.070 822.330 2076.970 822.390 ;
        RECT 2254.070 822.330 2256.970 822.390 ;
        RECT 2434.070 822.330 2436.970 822.390 ;
        RECT 2614.070 822.330 2616.970 822.390 ;
        RECT 2794.070 822.330 2796.970 822.390 ;
        RECT 2931.250 822.330 2934.150 822.390 ;
        RECT -14.530 819.430 2934.150 822.330 ;
        RECT -14.530 819.370 -11.630 819.430 ;
        RECT 94.070 819.370 96.970 819.430 ;
        RECT 274.070 819.370 276.970 819.430 ;
        RECT 454.070 819.370 456.970 819.430 ;
        RECT 634.070 819.370 636.970 819.430 ;
        RECT 814.070 819.370 816.970 819.430 ;
        RECT 994.070 819.370 996.970 819.430 ;
        RECT 1174.070 819.370 1176.970 819.430 ;
        RECT 1354.070 819.370 1356.970 819.430 ;
        RECT 1534.070 819.370 1536.970 819.430 ;
        RECT 1714.070 819.370 1716.970 819.430 ;
        RECT 1894.070 819.370 1896.970 819.430 ;
        RECT 2074.070 819.370 2076.970 819.430 ;
        RECT 2254.070 819.370 2256.970 819.430 ;
        RECT 2434.070 819.370 2436.970 819.430 ;
        RECT 2614.070 819.370 2616.970 819.430 ;
        RECT 2794.070 819.370 2796.970 819.430 ;
        RECT 2931.250 819.370 2934.150 819.430 ;
        RECT -14.530 642.330 -11.630 642.390 ;
        RECT 94.070 642.330 96.970 642.390 ;
        RECT 274.070 642.330 276.970 642.390 ;
        RECT 454.070 642.330 456.970 642.390 ;
        RECT 634.070 642.330 636.970 642.390 ;
        RECT 814.070 642.330 816.970 642.390 ;
        RECT 994.070 642.330 996.970 642.390 ;
        RECT 1174.070 642.330 1176.970 642.390 ;
        RECT 1354.070 642.330 1356.970 642.390 ;
        RECT 1534.070 642.330 1536.970 642.390 ;
        RECT 1714.070 642.330 1716.970 642.390 ;
        RECT 1894.070 642.330 1896.970 642.390 ;
        RECT 2074.070 642.330 2076.970 642.390 ;
        RECT 2254.070 642.330 2256.970 642.390 ;
        RECT 2434.070 642.330 2436.970 642.390 ;
        RECT 2614.070 642.330 2616.970 642.390 ;
        RECT 2794.070 642.330 2796.970 642.390 ;
        RECT 2931.250 642.330 2934.150 642.390 ;
        RECT -14.530 639.430 2934.150 642.330 ;
        RECT -14.530 639.370 -11.630 639.430 ;
        RECT 94.070 639.370 96.970 639.430 ;
        RECT 274.070 639.370 276.970 639.430 ;
        RECT 454.070 639.370 456.970 639.430 ;
        RECT 634.070 639.370 636.970 639.430 ;
        RECT 814.070 639.370 816.970 639.430 ;
        RECT 994.070 639.370 996.970 639.430 ;
        RECT 1174.070 639.370 1176.970 639.430 ;
        RECT 1354.070 639.370 1356.970 639.430 ;
        RECT 1534.070 639.370 1536.970 639.430 ;
        RECT 1714.070 639.370 1716.970 639.430 ;
        RECT 1894.070 639.370 1896.970 639.430 ;
        RECT 2074.070 639.370 2076.970 639.430 ;
        RECT 2254.070 639.370 2256.970 639.430 ;
        RECT 2434.070 639.370 2436.970 639.430 ;
        RECT 2614.070 639.370 2616.970 639.430 ;
        RECT 2794.070 639.370 2796.970 639.430 ;
        RECT 2931.250 639.370 2934.150 639.430 ;
        RECT -14.530 462.330 -11.630 462.390 ;
        RECT 94.070 462.330 96.970 462.390 ;
        RECT 274.070 462.330 276.970 462.390 ;
        RECT 454.070 462.330 456.970 462.390 ;
        RECT 634.070 462.330 636.970 462.390 ;
        RECT 814.070 462.330 816.970 462.390 ;
        RECT 994.070 462.330 996.970 462.390 ;
        RECT 1174.070 462.330 1176.970 462.390 ;
        RECT 1354.070 462.330 1356.970 462.390 ;
        RECT 1534.070 462.330 1536.970 462.390 ;
        RECT 1714.070 462.330 1716.970 462.390 ;
        RECT 1894.070 462.330 1896.970 462.390 ;
        RECT 2074.070 462.330 2076.970 462.390 ;
        RECT 2254.070 462.330 2256.970 462.390 ;
        RECT 2434.070 462.330 2436.970 462.390 ;
        RECT 2614.070 462.330 2616.970 462.390 ;
        RECT 2794.070 462.330 2796.970 462.390 ;
        RECT 2931.250 462.330 2934.150 462.390 ;
        RECT -14.530 459.430 2934.150 462.330 ;
        RECT -14.530 459.370 -11.630 459.430 ;
        RECT 94.070 459.370 96.970 459.430 ;
        RECT 274.070 459.370 276.970 459.430 ;
        RECT 454.070 459.370 456.970 459.430 ;
        RECT 634.070 459.370 636.970 459.430 ;
        RECT 814.070 459.370 816.970 459.430 ;
        RECT 994.070 459.370 996.970 459.430 ;
        RECT 1174.070 459.370 1176.970 459.430 ;
        RECT 1354.070 459.370 1356.970 459.430 ;
        RECT 1534.070 459.370 1536.970 459.430 ;
        RECT 1714.070 459.370 1716.970 459.430 ;
        RECT 1894.070 459.370 1896.970 459.430 ;
        RECT 2074.070 459.370 2076.970 459.430 ;
        RECT 2254.070 459.370 2256.970 459.430 ;
        RECT 2434.070 459.370 2436.970 459.430 ;
        RECT 2614.070 459.370 2616.970 459.430 ;
        RECT 2794.070 459.370 2796.970 459.430 ;
        RECT 2931.250 459.370 2934.150 459.430 ;
        RECT -14.530 282.330 -11.630 282.390 ;
        RECT 94.070 282.330 96.970 282.390 ;
        RECT 274.070 282.330 276.970 282.390 ;
        RECT 454.070 282.330 456.970 282.390 ;
        RECT 634.070 282.330 636.970 282.390 ;
        RECT 814.070 282.330 816.970 282.390 ;
        RECT 994.070 282.330 996.970 282.390 ;
        RECT 1174.070 282.330 1176.970 282.390 ;
        RECT 1354.070 282.330 1356.970 282.390 ;
        RECT 1534.070 282.330 1536.970 282.390 ;
        RECT 1714.070 282.330 1716.970 282.390 ;
        RECT 1894.070 282.330 1896.970 282.390 ;
        RECT 2074.070 282.330 2076.970 282.390 ;
        RECT 2254.070 282.330 2256.970 282.390 ;
        RECT 2434.070 282.330 2436.970 282.390 ;
        RECT 2614.070 282.330 2616.970 282.390 ;
        RECT 2794.070 282.330 2796.970 282.390 ;
        RECT 2931.250 282.330 2934.150 282.390 ;
        RECT -14.530 279.430 2934.150 282.330 ;
        RECT -14.530 279.370 -11.630 279.430 ;
        RECT 94.070 279.370 96.970 279.430 ;
        RECT 274.070 279.370 276.970 279.430 ;
        RECT 454.070 279.370 456.970 279.430 ;
        RECT 634.070 279.370 636.970 279.430 ;
        RECT 814.070 279.370 816.970 279.430 ;
        RECT 994.070 279.370 996.970 279.430 ;
        RECT 1174.070 279.370 1176.970 279.430 ;
        RECT 1354.070 279.370 1356.970 279.430 ;
        RECT 1534.070 279.370 1536.970 279.430 ;
        RECT 1714.070 279.370 1716.970 279.430 ;
        RECT 1894.070 279.370 1896.970 279.430 ;
        RECT 2074.070 279.370 2076.970 279.430 ;
        RECT 2254.070 279.370 2256.970 279.430 ;
        RECT 2434.070 279.370 2436.970 279.430 ;
        RECT 2614.070 279.370 2616.970 279.430 ;
        RECT 2794.070 279.370 2796.970 279.430 ;
        RECT 2931.250 279.370 2934.150 279.430 ;
        RECT -14.530 102.330 -11.630 102.390 ;
        RECT 94.070 102.330 96.970 102.390 ;
        RECT 274.070 102.330 276.970 102.390 ;
        RECT 454.070 102.330 456.970 102.390 ;
        RECT 634.070 102.330 636.970 102.390 ;
        RECT 814.070 102.330 816.970 102.390 ;
        RECT 994.070 102.330 996.970 102.390 ;
        RECT 1174.070 102.330 1176.970 102.390 ;
        RECT 1354.070 102.330 1356.970 102.390 ;
        RECT 1534.070 102.330 1536.970 102.390 ;
        RECT 1714.070 102.330 1716.970 102.390 ;
        RECT 1894.070 102.330 1896.970 102.390 ;
        RECT 2074.070 102.330 2076.970 102.390 ;
        RECT 2254.070 102.330 2256.970 102.390 ;
        RECT 2434.070 102.330 2436.970 102.390 ;
        RECT 2614.070 102.330 2616.970 102.390 ;
        RECT 2794.070 102.330 2796.970 102.390 ;
        RECT 2931.250 102.330 2934.150 102.390 ;
        RECT -14.530 99.430 2934.150 102.330 ;
        RECT -14.530 99.370 -11.630 99.430 ;
        RECT 94.070 99.370 96.970 99.430 ;
        RECT 274.070 99.370 276.970 99.430 ;
        RECT 454.070 99.370 456.970 99.430 ;
        RECT 634.070 99.370 636.970 99.430 ;
        RECT 814.070 99.370 816.970 99.430 ;
        RECT 994.070 99.370 996.970 99.430 ;
        RECT 1174.070 99.370 1176.970 99.430 ;
        RECT 1354.070 99.370 1356.970 99.430 ;
        RECT 1534.070 99.370 1536.970 99.430 ;
        RECT 1714.070 99.370 1716.970 99.430 ;
        RECT 1894.070 99.370 1896.970 99.430 ;
        RECT 2074.070 99.370 2076.970 99.430 ;
        RECT 2254.070 99.370 2256.970 99.430 ;
        RECT 2434.070 99.370 2436.970 99.430 ;
        RECT 2614.070 99.370 2616.970 99.430 ;
        RECT 2794.070 99.370 2796.970 99.430 ;
        RECT 2931.250 99.370 2934.150 99.430 ;
        RECT -14.530 -6.270 -11.630 -6.210 ;
        RECT 94.070 -6.270 96.970 -6.210 ;
        RECT 274.070 -6.270 276.970 -6.210 ;
        RECT 454.070 -6.270 456.970 -6.210 ;
        RECT 634.070 -6.270 636.970 -6.210 ;
        RECT 814.070 -6.270 816.970 -6.210 ;
        RECT 994.070 -6.270 996.970 -6.210 ;
        RECT 1174.070 -6.270 1176.970 -6.210 ;
        RECT 1354.070 -6.270 1356.970 -6.210 ;
        RECT 1534.070 -6.270 1536.970 -6.210 ;
        RECT 1714.070 -6.270 1716.970 -6.210 ;
        RECT 1894.070 -6.270 1896.970 -6.210 ;
        RECT 2074.070 -6.270 2076.970 -6.210 ;
        RECT 2254.070 -6.270 2256.970 -6.210 ;
        RECT 2434.070 -6.270 2436.970 -6.210 ;
        RECT 2614.070 -6.270 2616.970 -6.210 ;
        RECT 2794.070 -6.270 2796.970 -6.210 ;
        RECT 2931.250 -6.270 2934.150 -6.210 ;
        RECT -14.530 -9.170 2934.150 -6.270 ;
        RECT -14.530 -9.230 -11.630 -9.170 ;
        RECT 94.070 -9.230 96.970 -9.170 ;
        RECT 274.070 -9.230 276.970 -9.170 ;
        RECT 454.070 -9.230 456.970 -9.170 ;
        RECT 634.070 -9.230 636.970 -9.170 ;
        RECT 814.070 -9.230 816.970 -9.170 ;
        RECT 994.070 -9.230 996.970 -9.170 ;
        RECT 1174.070 -9.230 1176.970 -9.170 ;
        RECT 1354.070 -9.230 1356.970 -9.170 ;
        RECT 1534.070 -9.230 1536.970 -9.170 ;
        RECT 1714.070 -9.230 1716.970 -9.170 ;
        RECT 1894.070 -9.230 1896.970 -9.170 ;
        RECT 2074.070 -9.230 2076.970 -9.170 ;
        RECT 2254.070 -9.230 2256.970 -9.170 ;
        RECT 2434.070 -9.230 2436.970 -9.170 ;
        RECT 2614.070 -9.230 2616.970 -9.170 ;
        RECT 2794.070 -9.230 2796.970 -9.170 ;
        RECT 2931.250 -9.230 2934.150 -9.170 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.130 -13.770 -16.230 3533.450 ;
        RECT 21.470 -18.370 24.370 3538.050 ;
        RECT 201.470 -18.370 204.370 3538.050 ;
        RECT 381.470 -18.370 384.370 3538.050 ;
        RECT 561.470 -18.370 564.370 3538.050 ;
        RECT 741.470 -18.370 744.370 3538.050 ;
        RECT 921.470 -18.370 924.370 3538.050 ;
        RECT 1101.470 -18.370 1104.370 3538.050 ;
        RECT 1281.470 -18.370 1284.370 3538.050 ;
        RECT 1461.470 -18.370 1464.370 3538.050 ;
        RECT 1641.470 -18.370 1644.370 3538.050 ;
        RECT 1821.470 -18.370 1824.370 3538.050 ;
        RECT 2001.470 -18.370 2004.370 3538.050 ;
        RECT 2181.470 -18.370 2184.370 3538.050 ;
        RECT 2361.470 -18.370 2364.370 3538.050 ;
        RECT 2541.470 -18.370 2544.370 3538.050 ;
        RECT 2721.470 -18.370 2724.370 3538.050 ;
        RECT 2901.470 -18.370 2904.370 3538.050 ;
        RECT 2935.850 -13.770 2938.750 3533.450 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3448.490 -17.090 3449.670 ;
        RECT -18.270 3446.890 -17.090 3448.070 ;
        RECT -18.270 3268.490 -17.090 3269.670 ;
        RECT -18.270 3266.890 -17.090 3268.070 ;
        RECT -18.270 3088.490 -17.090 3089.670 ;
        RECT -18.270 3086.890 -17.090 3088.070 ;
        RECT -18.270 2908.490 -17.090 2909.670 ;
        RECT -18.270 2906.890 -17.090 2908.070 ;
        RECT -18.270 2728.490 -17.090 2729.670 ;
        RECT -18.270 2726.890 -17.090 2728.070 ;
        RECT -18.270 2548.490 -17.090 2549.670 ;
        RECT -18.270 2546.890 -17.090 2548.070 ;
        RECT -18.270 2368.490 -17.090 2369.670 ;
        RECT -18.270 2366.890 -17.090 2368.070 ;
        RECT -18.270 2188.490 -17.090 2189.670 ;
        RECT -18.270 2186.890 -17.090 2188.070 ;
        RECT -18.270 2008.490 -17.090 2009.670 ;
        RECT -18.270 2006.890 -17.090 2008.070 ;
        RECT -18.270 1828.490 -17.090 1829.670 ;
        RECT -18.270 1826.890 -17.090 1828.070 ;
        RECT -18.270 1648.490 -17.090 1649.670 ;
        RECT -18.270 1646.890 -17.090 1648.070 ;
        RECT -18.270 1468.490 -17.090 1469.670 ;
        RECT -18.270 1466.890 -17.090 1468.070 ;
        RECT -18.270 1288.490 -17.090 1289.670 ;
        RECT -18.270 1286.890 -17.090 1288.070 ;
        RECT -18.270 1108.490 -17.090 1109.670 ;
        RECT -18.270 1106.890 -17.090 1108.070 ;
        RECT -18.270 928.490 -17.090 929.670 ;
        RECT -18.270 926.890 -17.090 928.070 ;
        RECT -18.270 748.490 -17.090 749.670 ;
        RECT -18.270 746.890 -17.090 748.070 ;
        RECT -18.270 568.490 -17.090 569.670 ;
        RECT -18.270 566.890 -17.090 568.070 ;
        RECT -18.270 388.490 -17.090 389.670 ;
        RECT -18.270 386.890 -17.090 388.070 ;
        RECT -18.270 208.490 -17.090 209.670 ;
        RECT -18.270 206.890 -17.090 208.070 ;
        RECT -18.270 28.490 -17.090 29.670 ;
        RECT -18.270 26.890 -17.090 28.070 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.330 3532.210 23.510 3533.390 ;
        RECT 22.330 3530.610 23.510 3531.790 ;
        RECT 22.330 3448.490 23.510 3449.670 ;
        RECT 22.330 3446.890 23.510 3448.070 ;
        RECT 22.330 3268.490 23.510 3269.670 ;
        RECT 22.330 3266.890 23.510 3268.070 ;
        RECT 22.330 3088.490 23.510 3089.670 ;
        RECT 22.330 3086.890 23.510 3088.070 ;
        RECT 22.330 2908.490 23.510 2909.670 ;
        RECT 22.330 2906.890 23.510 2908.070 ;
        RECT 22.330 2728.490 23.510 2729.670 ;
        RECT 22.330 2726.890 23.510 2728.070 ;
        RECT 22.330 2548.490 23.510 2549.670 ;
        RECT 22.330 2546.890 23.510 2548.070 ;
        RECT 22.330 2368.490 23.510 2369.670 ;
        RECT 22.330 2366.890 23.510 2368.070 ;
        RECT 22.330 2188.490 23.510 2189.670 ;
        RECT 22.330 2186.890 23.510 2188.070 ;
        RECT 22.330 2008.490 23.510 2009.670 ;
        RECT 22.330 2006.890 23.510 2008.070 ;
        RECT 22.330 1828.490 23.510 1829.670 ;
        RECT 22.330 1826.890 23.510 1828.070 ;
        RECT 22.330 1648.490 23.510 1649.670 ;
        RECT 22.330 1646.890 23.510 1648.070 ;
        RECT 22.330 1468.490 23.510 1469.670 ;
        RECT 22.330 1466.890 23.510 1468.070 ;
        RECT 22.330 1288.490 23.510 1289.670 ;
        RECT 22.330 1286.890 23.510 1288.070 ;
        RECT 22.330 1108.490 23.510 1109.670 ;
        RECT 22.330 1106.890 23.510 1108.070 ;
        RECT 22.330 928.490 23.510 929.670 ;
        RECT 22.330 926.890 23.510 928.070 ;
        RECT 22.330 748.490 23.510 749.670 ;
        RECT 22.330 746.890 23.510 748.070 ;
        RECT 22.330 568.490 23.510 569.670 ;
        RECT 22.330 566.890 23.510 568.070 ;
        RECT 22.330 388.490 23.510 389.670 ;
        RECT 22.330 386.890 23.510 388.070 ;
        RECT 22.330 208.490 23.510 209.670 ;
        RECT 22.330 206.890 23.510 208.070 ;
        RECT 22.330 28.490 23.510 29.670 ;
        RECT 22.330 26.890 23.510 28.070 ;
        RECT 22.330 -12.110 23.510 -10.930 ;
        RECT 22.330 -13.710 23.510 -12.530 ;
        RECT 202.330 3532.210 203.510 3533.390 ;
        RECT 202.330 3530.610 203.510 3531.790 ;
        RECT 202.330 3448.490 203.510 3449.670 ;
        RECT 202.330 3446.890 203.510 3448.070 ;
        RECT 202.330 3268.490 203.510 3269.670 ;
        RECT 202.330 3266.890 203.510 3268.070 ;
        RECT 202.330 3088.490 203.510 3089.670 ;
        RECT 202.330 3086.890 203.510 3088.070 ;
        RECT 202.330 2908.490 203.510 2909.670 ;
        RECT 202.330 2906.890 203.510 2908.070 ;
        RECT 202.330 2728.490 203.510 2729.670 ;
        RECT 202.330 2726.890 203.510 2728.070 ;
        RECT 202.330 2548.490 203.510 2549.670 ;
        RECT 202.330 2546.890 203.510 2548.070 ;
        RECT 202.330 2368.490 203.510 2369.670 ;
        RECT 202.330 2366.890 203.510 2368.070 ;
        RECT 202.330 2188.490 203.510 2189.670 ;
        RECT 202.330 2186.890 203.510 2188.070 ;
        RECT 202.330 2008.490 203.510 2009.670 ;
        RECT 202.330 2006.890 203.510 2008.070 ;
        RECT 202.330 1828.490 203.510 1829.670 ;
        RECT 202.330 1826.890 203.510 1828.070 ;
        RECT 202.330 1648.490 203.510 1649.670 ;
        RECT 202.330 1646.890 203.510 1648.070 ;
        RECT 202.330 1468.490 203.510 1469.670 ;
        RECT 202.330 1466.890 203.510 1468.070 ;
        RECT 202.330 1288.490 203.510 1289.670 ;
        RECT 202.330 1286.890 203.510 1288.070 ;
        RECT 202.330 1108.490 203.510 1109.670 ;
        RECT 202.330 1106.890 203.510 1108.070 ;
        RECT 202.330 928.490 203.510 929.670 ;
        RECT 202.330 926.890 203.510 928.070 ;
        RECT 202.330 748.490 203.510 749.670 ;
        RECT 202.330 746.890 203.510 748.070 ;
        RECT 202.330 568.490 203.510 569.670 ;
        RECT 202.330 566.890 203.510 568.070 ;
        RECT 202.330 388.490 203.510 389.670 ;
        RECT 202.330 386.890 203.510 388.070 ;
        RECT 202.330 208.490 203.510 209.670 ;
        RECT 202.330 206.890 203.510 208.070 ;
        RECT 202.330 28.490 203.510 29.670 ;
        RECT 202.330 26.890 203.510 28.070 ;
        RECT 202.330 -12.110 203.510 -10.930 ;
        RECT 202.330 -13.710 203.510 -12.530 ;
        RECT 382.330 3532.210 383.510 3533.390 ;
        RECT 382.330 3530.610 383.510 3531.790 ;
        RECT 382.330 3448.490 383.510 3449.670 ;
        RECT 382.330 3446.890 383.510 3448.070 ;
        RECT 382.330 3268.490 383.510 3269.670 ;
        RECT 382.330 3266.890 383.510 3268.070 ;
        RECT 382.330 3088.490 383.510 3089.670 ;
        RECT 382.330 3086.890 383.510 3088.070 ;
        RECT 382.330 2908.490 383.510 2909.670 ;
        RECT 382.330 2906.890 383.510 2908.070 ;
        RECT 382.330 2728.490 383.510 2729.670 ;
        RECT 382.330 2726.890 383.510 2728.070 ;
        RECT 382.330 2548.490 383.510 2549.670 ;
        RECT 382.330 2546.890 383.510 2548.070 ;
        RECT 382.330 2368.490 383.510 2369.670 ;
        RECT 382.330 2366.890 383.510 2368.070 ;
        RECT 382.330 2188.490 383.510 2189.670 ;
        RECT 382.330 2186.890 383.510 2188.070 ;
        RECT 382.330 2008.490 383.510 2009.670 ;
        RECT 382.330 2006.890 383.510 2008.070 ;
        RECT 382.330 1828.490 383.510 1829.670 ;
        RECT 382.330 1826.890 383.510 1828.070 ;
        RECT 382.330 1648.490 383.510 1649.670 ;
        RECT 382.330 1646.890 383.510 1648.070 ;
        RECT 382.330 1468.490 383.510 1469.670 ;
        RECT 382.330 1466.890 383.510 1468.070 ;
        RECT 382.330 1288.490 383.510 1289.670 ;
        RECT 382.330 1286.890 383.510 1288.070 ;
        RECT 382.330 1108.490 383.510 1109.670 ;
        RECT 382.330 1106.890 383.510 1108.070 ;
        RECT 382.330 928.490 383.510 929.670 ;
        RECT 382.330 926.890 383.510 928.070 ;
        RECT 382.330 748.490 383.510 749.670 ;
        RECT 382.330 746.890 383.510 748.070 ;
        RECT 382.330 568.490 383.510 569.670 ;
        RECT 382.330 566.890 383.510 568.070 ;
        RECT 382.330 388.490 383.510 389.670 ;
        RECT 382.330 386.890 383.510 388.070 ;
        RECT 382.330 208.490 383.510 209.670 ;
        RECT 382.330 206.890 383.510 208.070 ;
        RECT 382.330 28.490 383.510 29.670 ;
        RECT 382.330 26.890 383.510 28.070 ;
        RECT 382.330 -12.110 383.510 -10.930 ;
        RECT 382.330 -13.710 383.510 -12.530 ;
        RECT 562.330 3532.210 563.510 3533.390 ;
        RECT 562.330 3530.610 563.510 3531.790 ;
        RECT 562.330 3448.490 563.510 3449.670 ;
        RECT 562.330 3446.890 563.510 3448.070 ;
        RECT 562.330 3268.490 563.510 3269.670 ;
        RECT 562.330 3266.890 563.510 3268.070 ;
        RECT 562.330 3088.490 563.510 3089.670 ;
        RECT 562.330 3086.890 563.510 3088.070 ;
        RECT 562.330 2908.490 563.510 2909.670 ;
        RECT 562.330 2906.890 563.510 2908.070 ;
        RECT 562.330 2728.490 563.510 2729.670 ;
        RECT 562.330 2726.890 563.510 2728.070 ;
        RECT 562.330 2548.490 563.510 2549.670 ;
        RECT 562.330 2546.890 563.510 2548.070 ;
        RECT 562.330 2368.490 563.510 2369.670 ;
        RECT 562.330 2366.890 563.510 2368.070 ;
        RECT 562.330 2188.490 563.510 2189.670 ;
        RECT 562.330 2186.890 563.510 2188.070 ;
        RECT 562.330 2008.490 563.510 2009.670 ;
        RECT 562.330 2006.890 563.510 2008.070 ;
        RECT 562.330 1828.490 563.510 1829.670 ;
        RECT 562.330 1826.890 563.510 1828.070 ;
        RECT 562.330 1648.490 563.510 1649.670 ;
        RECT 562.330 1646.890 563.510 1648.070 ;
        RECT 562.330 1468.490 563.510 1469.670 ;
        RECT 562.330 1466.890 563.510 1468.070 ;
        RECT 562.330 1288.490 563.510 1289.670 ;
        RECT 562.330 1286.890 563.510 1288.070 ;
        RECT 562.330 1108.490 563.510 1109.670 ;
        RECT 562.330 1106.890 563.510 1108.070 ;
        RECT 562.330 928.490 563.510 929.670 ;
        RECT 562.330 926.890 563.510 928.070 ;
        RECT 562.330 748.490 563.510 749.670 ;
        RECT 562.330 746.890 563.510 748.070 ;
        RECT 562.330 568.490 563.510 569.670 ;
        RECT 562.330 566.890 563.510 568.070 ;
        RECT 562.330 388.490 563.510 389.670 ;
        RECT 562.330 386.890 563.510 388.070 ;
        RECT 562.330 208.490 563.510 209.670 ;
        RECT 562.330 206.890 563.510 208.070 ;
        RECT 562.330 28.490 563.510 29.670 ;
        RECT 562.330 26.890 563.510 28.070 ;
        RECT 562.330 -12.110 563.510 -10.930 ;
        RECT 562.330 -13.710 563.510 -12.530 ;
        RECT 742.330 3532.210 743.510 3533.390 ;
        RECT 742.330 3530.610 743.510 3531.790 ;
        RECT 742.330 3448.490 743.510 3449.670 ;
        RECT 742.330 3446.890 743.510 3448.070 ;
        RECT 742.330 3268.490 743.510 3269.670 ;
        RECT 742.330 3266.890 743.510 3268.070 ;
        RECT 742.330 3088.490 743.510 3089.670 ;
        RECT 742.330 3086.890 743.510 3088.070 ;
        RECT 742.330 2908.490 743.510 2909.670 ;
        RECT 742.330 2906.890 743.510 2908.070 ;
        RECT 742.330 2728.490 743.510 2729.670 ;
        RECT 742.330 2726.890 743.510 2728.070 ;
        RECT 742.330 2548.490 743.510 2549.670 ;
        RECT 742.330 2546.890 743.510 2548.070 ;
        RECT 742.330 2368.490 743.510 2369.670 ;
        RECT 742.330 2366.890 743.510 2368.070 ;
        RECT 742.330 2188.490 743.510 2189.670 ;
        RECT 742.330 2186.890 743.510 2188.070 ;
        RECT 742.330 2008.490 743.510 2009.670 ;
        RECT 742.330 2006.890 743.510 2008.070 ;
        RECT 742.330 1828.490 743.510 1829.670 ;
        RECT 742.330 1826.890 743.510 1828.070 ;
        RECT 742.330 1648.490 743.510 1649.670 ;
        RECT 742.330 1646.890 743.510 1648.070 ;
        RECT 742.330 1468.490 743.510 1469.670 ;
        RECT 742.330 1466.890 743.510 1468.070 ;
        RECT 742.330 1288.490 743.510 1289.670 ;
        RECT 742.330 1286.890 743.510 1288.070 ;
        RECT 742.330 1108.490 743.510 1109.670 ;
        RECT 742.330 1106.890 743.510 1108.070 ;
        RECT 742.330 928.490 743.510 929.670 ;
        RECT 742.330 926.890 743.510 928.070 ;
        RECT 742.330 748.490 743.510 749.670 ;
        RECT 742.330 746.890 743.510 748.070 ;
        RECT 742.330 568.490 743.510 569.670 ;
        RECT 742.330 566.890 743.510 568.070 ;
        RECT 742.330 388.490 743.510 389.670 ;
        RECT 742.330 386.890 743.510 388.070 ;
        RECT 742.330 208.490 743.510 209.670 ;
        RECT 742.330 206.890 743.510 208.070 ;
        RECT 742.330 28.490 743.510 29.670 ;
        RECT 742.330 26.890 743.510 28.070 ;
        RECT 742.330 -12.110 743.510 -10.930 ;
        RECT 742.330 -13.710 743.510 -12.530 ;
        RECT 922.330 3532.210 923.510 3533.390 ;
        RECT 922.330 3530.610 923.510 3531.790 ;
        RECT 922.330 3448.490 923.510 3449.670 ;
        RECT 922.330 3446.890 923.510 3448.070 ;
        RECT 922.330 3268.490 923.510 3269.670 ;
        RECT 922.330 3266.890 923.510 3268.070 ;
        RECT 922.330 3088.490 923.510 3089.670 ;
        RECT 922.330 3086.890 923.510 3088.070 ;
        RECT 922.330 2908.490 923.510 2909.670 ;
        RECT 922.330 2906.890 923.510 2908.070 ;
        RECT 922.330 2728.490 923.510 2729.670 ;
        RECT 922.330 2726.890 923.510 2728.070 ;
        RECT 922.330 2548.490 923.510 2549.670 ;
        RECT 922.330 2546.890 923.510 2548.070 ;
        RECT 922.330 2368.490 923.510 2369.670 ;
        RECT 922.330 2366.890 923.510 2368.070 ;
        RECT 922.330 2188.490 923.510 2189.670 ;
        RECT 922.330 2186.890 923.510 2188.070 ;
        RECT 922.330 2008.490 923.510 2009.670 ;
        RECT 922.330 2006.890 923.510 2008.070 ;
        RECT 922.330 1828.490 923.510 1829.670 ;
        RECT 922.330 1826.890 923.510 1828.070 ;
        RECT 922.330 1648.490 923.510 1649.670 ;
        RECT 922.330 1646.890 923.510 1648.070 ;
        RECT 922.330 1468.490 923.510 1469.670 ;
        RECT 922.330 1466.890 923.510 1468.070 ;
        RECT 922.330 1288.490 923.510 1289.670 ;
        RECT 922.330 1286.890 923.510 1288.070 ;
        RECT 922.330 1108.490 923.510 1109.670 ;
        RECT 922.330 1106.890 923.510 1108.070 ;
        RECT 922.330 928.490 923.510 929.670 ;
        RECT 922.330 926.890 923.510 928.070 ;
        RECT 922.330 748.490 923.510 749.670 ;
        RECT 922.330 746.890 923.510 748.070 ;
        RECT 922.330 568.490 923.510 569.670 ;
        RECT 922.330 566.890 923.510 568.070 ;
        RECT 922.330 388.490 923.510 389.670 ;
        RECT 922.330 386.890 923.510 388.070 ;
        RECT 922.330 208.490 923.510 209.670 ;
        RECT 922.330 206.890 923.510 208.070 ;
        RECT 922.330 28.490 923.510 29.670 ;
        RECT 922.330 26.890 923.510 28.070 ;
        RECT 922.330 -12.110 923.510 -10.930 ;
        RECT 922.330 -13.710 923.510 -12.530 ;
        RECT 1102.330 3532.210 1103.510 3533.390 ;
        RECT 1102.330 3530.610 1103.510 3531.790 ;
        RECT 1102.330 3448.490 1103.510 3449.670 ;
        RECT 1102.330 3446.890 1103.510 3448.070 ;
        RECT 1102.330 3268.490 1103.510 3269.670 ;
        RECT 1102.330 3266.890 1103.510 3268.070 ;
        RECT 1102.330 3088.490 1103.510 3089.670 ;
        RECT 1102.330 3086.890 1103.510 3088.070 ;
        RECT 1102.330 2908.490 1103.510 2909.670 ;
        RECT 1102.330 2906.890 1103.510 2908.070 ;
        RECT 1102.330 2728.490 1103.510 2729.670 ;
        RECT 1102.330 2726.890 1103.510 2728.070 ;
        RECT 1102.330 2548.490 1103.510 2549.670 ;
        RECT 1102.330 2546.890 1103.510 2548.070 ;
        RECT 1102.330 2368.490 1103.510 2369.670 ;
        RECT 1102.330 2366.890 1103.510 2368.070 ;
        RECT 1102.330 2188.490 1103.510 2189.670 ;
        RECT 1102.330 2186.890 1103.510 2188.070 ;
        RECT 1102.330 2008.490 1103.510 2009.670 ;
        RECT 1102.330 2006.890 1103.510 2008.070 ;
        RECT 1102.330 1828.490 1103.510 1829.670 ;
        RECT 1102.330 1826.890 1103.510 1828.070 ;
        RECT 1102.330 1648.490 1103.510 1649.670 ;
        RECT 1102.330 1646.890 1103.510 1648.070 ;
        RECT 1102.330 1468.490 1103.510 1469.670 ;
        RECT 1102.330 1466.890 1103.510 1468.070 ;
        RECT 1102.330 1288.490 1103.510 1289.670 ;
        RECT 1102.330 1286.890 1103.510 1288.070 ;
        RECT 1102.330 1108.490 1103.510 1109.670 ;
        RECT 1102.330 1106.890 1103.510 1108.070 ;
        RECT 1102.330 928.490 1103.510 929.670 ;
        RECT 1102.330 926.890 1103.510 928.070 ;
        RECT 1102.330 748.490 1103.510 749.670 ;
        RECT 1102.330 746.890 1103.510 748.070 ;
        RECT 1102.330 568.490 1103.510 569.670 ;
        RECT 1102.330 566.890 1103.510 568.070 ;
        RECT 1102.330 388.490 1103.510 389.670 ;
        RECT 1102.330 386.890 1103.510 388.070 ;
        RECT 1102.330 208.490 1103.510 209.670 ;
        RECT 1102.330 206.890 1103.510 208.070 ;
        RECT 1102.330 28.490 1103.510 29.670 ;
        RECT 1102.330 26.890 1103.510 28.070 ;
        RECT 1102.330 -12.110 1103.510 -10.930 ;
        RECT 1102.330 -13.710 1103.510 -12.530 ;
        RECT 1282.330 3532.210 1283.510 3533.390 ;
        RECT 1282.330 3530.610 1283.510 3531.790 ;
        RECT 1282.330 3448.490 1283.510 3449.670 ;
        RECT 1282.330 3446.890 1283.510 3448.070 ;
        RECT 1282.330 3268.490 1283.510 3269.670 ;
        RECT 1282.330 3266.890 1283.510 3268.070 ;
        RECT 1282.330 3088.490 1283.510 3089.670 ;
        RECT 1282.330 3086.890 1283.510 3088.070 ;
        RECT 1282.330 2908.490 1283.510 2909.670 ;
        RECT 1282.330 2906.890 1283.510 2908.070 ;
        RECT 1282.330 2728.490 1283.510 2729.670 ;
        RECT 1282.330 2726.890 1283.510 2728.070 ;
        RECT 1282.330 2548.490 1283.510 2549.670 ;
        RECT 1282.330 2546.890 1283.510 2548.070 ;
        RECT 1282.330 2368.490 1283.510 2369.670 ;
        RECT 1282.330 2366.890 1283.510 2368.070 ;
        RECT 1282.330 2188.490 1283.510 2189.670 ;
        RECT 1282.330 2186.890 1283.510 2188.070 ;
        RECT 1282.330 2008.490 1283.510 2009.670 ;
        RECT 1282.330 2006.890 1283.510 2008.070 ;
        RECT 1282.330 1828.490 1283.510 1829.670 ;
        RECT 1282.330 1826.890 1283.510 1828.070 ;
        RECT 1282.330 1648.490 1283.510 1649.670 ;
        RECT 1282.330 1646.890 1283.510 1648.070 ;
        RECT 1282.330 1468.490 1283.510 1469.670 ;
        RECT 1282.330 1466.890 1283.510 1468.070 ;
        RECT 1282.330 1288.490 1283.510 1289.670 ;
        RECT 1282.330 1286.890 1283.510 1288.070 ;
        RECT 1282.330 1108.490 1283.510 1109.670 ;
        RECT 1282.330 1106.890 1283.510 1108.070 ;
        RECT 1282.330 928.490 1283.510 929.670 ;
        RECT 1282.330 926.890 1283.510 928.070 ;
        RECT 1282.330 748.490 1283.510 749.670 ;
        RECT 1282.330 746.890 1283.510 748.070 ;
        RECT 1282.330 568.490 1283.510 569.670 ;
        RECT 1282.330 566.890 1283.510 568.070 ;
        RECT 1282.330 388.490 1283.510 389.670 ;
        RECT 1282.330 386.890 1283.510 388.070 ;
        RECT 1282.330 208.490 1283.510 209.670 ;
        RECT 1282.330 206.890 1283.510 208.070 ;
        RECT 1282.330 28.490 1283.510 29.670 ;
        RECT 1282.330 26.890 1283.510 28.070 ;
        RECT 1282.330 -12.110 1283.510 -10.930 ;
        RECT 1282.330 -13.710 1283.510 -12.530 ;
        RECT 1462.330 3532.210 1463.510 3533.390 ;
        RECT 1462.330 3530.610 1463.510 3531.790 ;
        RECT 1462.330 3448.490 1463.510 3449.670 ;
        RECT 1462.330 3446.890 1463.510 3448.070 ;
        RECT 1462.330 3268.490 1463.510 3269.670 ;
        RECT 1462.330 3266.890 1463.510 3268.070 ;
        RECT 1462.330 3088.490 1463.510 3089.670 ;
        RECT 1462.330 3086.890 1463.510 3088.070 ;
        RECT 1462.330 2908.490 1463.510 2909.670 ;
        RECT 1462.330 2906.890 1463.510 2908.070 ;
        RECT 1462.330 2728.490 1463.510 2729.670 ;
        RECT 1462.330 2726.890 1463.510 2728.070 ;
        RECT 1462.330 2548.490 1463.510 2549.670 ;
        RECT 1462.330 2546.890 1463.510 2548.070 ;
        RECT 1462.330 2368.490 1463.510 2369.670 ;
        RECT 1462.330 2366.890 1463.510 2368.070 ;
        RECT 1462.330 2188.490 1463.510 2189.670 ;
        RECT 1462.330 2186.890 1463.510 2188.070 ;
        RECT 1462.330 2008.490 1463.510 2009.670 ;
        RECT 1462.330 2006.890 1463.510 2008.070 ;
        RECT 1462.330 1828.490 1463.510 1829.670 ;
        RECT 1462.330 1826.890 1463.510 1828.070 ;
        RECT 1462.330 1648.490 1463.510 1649.670 ;
        RECT 1462.330 1646.890 1463.510 1648.070 ;
        RECT 1462.330 1468.490 1463.510 1469.670 ;
        RECT 1462.330 1466.890 1463.510 1468.070 ;
        RECT 1462.330 1288.490 1463.510 1289.670 ;
        RECT 1462.330 1286.890 1463.510 1288.070 ;
        RECT 1462.330 1108.490 1463.510 1109.670 ;
        RECT 1462.330 1106.890 1463.510 1108.070 ;
        RECT 1462.330 928.490 1463.510 929.670 ;
        RECT 1462.330 926.890 1463.510 928.070 ;
        RECT 1462.330 748.490 1463.510 749.670 ;
        RECT 1462.330 746.890 1463.510 748.070 ;
        RECT 1462.330 568.490 1463.510 569.670 ;
        RECT 1462.330 566.890 1463.510 568.070 ;
        RECT 1462.330 388.490 1463.510 389.670 ;
        RECT 1462.330 386.890 1463.510 388.070 ;
        RECT 1462.330 208.490 1463.510 209.670 ;
        RECT 1462.330 206.890 1463.510 208.070 ;
        RECT 1462.330 28.490 1463.510 29.670 ;
        RECT 1462.330 26.890 1463.510 28.070 ;
        RECT 1462.330 -12.110 1463.510 -10.930 ;
        RECT 1462.330 -13.710 1463.510 -12.530 ;
        RECT 1642.330 3532.210 1643.510 3533.390 ;
        RECT 1642.330 3530.610 1643.510 3531.790 ;
        RECT 1642.330 3448.490 1643.510 3449.670 ;
        RECT 1642.330 3446.890 1643.510 3448.070 ;
        RECT 1642.330 3268.490 1643.510 3269.670 ;
        RECT 1642.330 3266.890 1643.510 3268.070 ;
        RECT 1642.330 3088.490 1643.510 3089.670 ;
        RECT 1642.330 3086.890 1643.510 3088.070 ;
        RECT 1642.330 2908.490 1643.510 2909.670 ;
        RECT 1642.330 2906.890 1643.510 2908.070 ;
        RECT 1642.330 2728.490 1643.510 2729.670 ;
        RECT 1642.330 2726.890 1643.510 2728.070 ;
        RECT 1642.330 2548.490 1643.510 2549.670 ;
        RECT 1642.330 2546.890 1643.510 2548.070 ;
        RECT 1642.330 2368.490 1643.510 2369.670 ;
        RECT 1642.330 2366.890 1643.510 2368.070 ;
        RECT 1642.330 2188.490 1643.510 2189.670 ;
        RECT 1642.330 2186.890 1643.510 2188.070 ;
        RECT 1642.330 2008.490 1643.510 2009.670 ;
        RECT 1642.330 2006.890 1643.510 2008.070 ;
        RECT 1642.330 1828.490 1643.510 1829.670 ;
        RECT 1642.330 1826.890 1643.510 1828.070 ;
        RECT 1642.330 1648.490 1643.510 1649.670 ;
        RECT 1642.330 1646.890 1643.510 1648.070 ;
        RECT 1642.330 1468.490 1643.510 1469.670 ;
        RECT 1642.330 1466.890 1643.510 1468.070 ;
        RECT 1642.330 1288.490 1643.510 1289.670 ;
        RECT 1642.330 1286.890 1643.510 1288.070 ;
        RECT 1642.330 1108.490 1643.510 1109.670 ;
        RECT 1642.330 1106.890 1643.510 1108.070 ;
        RECT 1642.330 928.490 1643.510 929.670 ;
        RECT 1642.330 926.890 1643.510 928.070 ;
        RECT 1642.330 748.490 1643.510 749.670 ;
        RECT 1642.330 746.890 1643.510 748.070 ;
        RECT 1642.330 568.490 1643.510 569.670 ;
        RECT 1642.330 566.890 1643.510 568.070 ;
        RECT 1642.330 388.490 1643.510 389.670 ;
        RECT 1642.330 386.890 1643.510 388.070 ;
        RECT 1642.330 208.490 1643.510 209.670 ;
        RECT 1642.330 206.890 1643.510 208.070 ;
        RECT 1642.330 28.490 1643.510 29.670 ;
        RECT 1642.330 26.890 1643.510 28.070 ;
        RECT 1642.330 -12.110 1643.510 -10.930 ;
        RECT 1642.330 -13.710 1643.510 -12.530 ;
        RECT 1822.330 3532.210 1823.510 3533.390 ;
        RECT 1822.330 3530.610 1823.510 3531.790 ;
        RECT 1822.330 3448.490 1823.510 3449.670 ;
        RECT 1822.330 3446.890 1823.510 3448.070 ;
        RECT 1822.330 3268.490 1823.510 3269.670 ;
        RECT 1822.330 3266.890 1823.510 3268.070 ;
        RECT 1822.330 3088.490 1823.510 3089.670 ;
        RECT 1822.330 3086.890 1823.510 3088.070 ;
        RECT 1822.330 2908.490 1823.510 2909.670 ;
        RECT 1822.330 2906.890 1823.510 2908.070 ;
        RECT 1822.330 2728.490 1823.510 2729.670 ;
        RECT 1822.330 2726.890 1823.510 2728.070 ;
        RECT 1822.330 2548.490 1823.510 2549.670 ;
        RECT 1822.330 2546.890 1823.510 2548.070 ;
        RECT 1822.330 2368.490 1823.510 2369.670 ;
        RECT 1822.330 2366.890 1823.510 2368.070 ;
        RECT 1822.330 2188.490 1823.510 2189.670 ;
        RECT 1822.330 2186.890 1823.510 2188.070 ;
        RECT 1822.330 2008.490 1823.510 2009.670 ;
        RECT 1822.330 2006.890 1823.510 2008.070 ;
        RECT 1822.330 1828.490 1823.510 1829.670 ;
        RECT 1822.330 1826.890 1823.510 1828.070 ;
        RECT 1822.330 1648.490 1823.510 1649.670 ;
        RECT 1822.330 1646.890 1823.510 1648.070 ;
        RECT 1822.330 1468.490 1823.510 1469.670 ;
        RECT 1822.330 1466.890 1823.510 1468.070 ;
        RECT 1822.330 1288.490 1823.510 1289.670 ;
        RECT 1822.330 1286.890 1823.510 1288.070 ;
        RECT 1822.330 1108.490 1823.510 1109.670 ;
        RECT 1822.330 1106.890 1823.510 1108.070 ;
        RECT 1822.330 928.490 1823.510 929.670 ;
        RECT 1822.330 926.890 1823.510 928.070 ;
        RECT 1822.330 748.490 1823.510 749.670 ;
        RECT 1822.330 746.890 1823.510 748.070 ;
        RECT 1822.330 568.490 1823.510 569.670 ;
        RECT 1822.330 566.890 1823.510 568.070 ;
        RECT 1822.330 388.490 1823.510 389.670 ;
        RECT 1822.330 386.890 1823.510 388.070 ;
        RECT 1822.330 208.490 1823.510 209.670 ;
        RECT 1822.330 206.890 1823.510 208.070 ;
        RECT 1822.330 28.490 1823.510 29.670 ;
        RECT 1822.330 26.890 1823.510 28.070 ;
        RECT 1822.330 -12.110 1823.510 -10.930 ;
        RECT 1822.330 -13.710 1823.510 -12.530 ;
        RECT 2002.330 3532.210 2003.510 3533.390 ;
        RECT 2002.330 3530.610 2003.510 3531.790 ;
        RECT 2002.330 3448.490 2003.510 3449.670 ;
        RECT 2002.330 3446.890 2003.510 3448.070 ;
        RECT 2002.330 3268.490 2003.510 3269.670 ;
        RECT 2002.330 3266.890 2003.510 3268.070 ;
        RECT 2002.330 3088.490 2003.510 3089.670 ;
        RECT 2002.330 3086.890 2003.510 3088.070 ;
        RECT 2002.330 2908.490 2003.510 2909.670 ;
        RECT 2002.330 2906.890 2003.510 2908.070 ;
        RECT 2002.330 2728.490 2003.510 2729.670 ;
        RECT 2002.330 2726.890 2003.510 2728.070 ;
        RECT 2002.330 2548.490 2003.510 2549.670 ;
        RECT 2002.330 2546.890 2003.510 2548.070 ;
        RECT 2002.330 2368.490 2003.510 2369.670 ;
        RECT 2002.330 2366.890 2003.510 2368.070 ;
        RECT 2002.330 2188.490 2003.510 2189.670 ;
        RECT 2002.330 2186.890 2003.510 2188.070 ;
        RECT 2002.330 2008.490 2003.510 2009.670 ;
        RECT 2002.330 2006.890 2003.510 2008.070 ;
        RECT 2002.330 1828.490 2003.510 1829.670 ;
        RECT 2002.330 1826.890 2003.510 1828.070 ;
        RECT 2002.330 1648.490 2003.510 1649.670 ;
        RECT 2002.330 1646.890 2003.510 1648.070 ;
        RECT 2002.330 1468.490 2003.510 1469.670 ;
        RECT 2002.330 1466.890 2003.510 1468.070 ;
        RECT 2002.330 1288.490 2003.510 1289.670 ;
        RECT 2002.330 1286.890 2003.510 1288.070 ;
        RECT 2002.330 1108.490 2003.510 1109.670 ;
        RECT 2002.330 1106.890 2003.510 1108.070 ;
        RECT 2002.330 928.490 2003.510 929.670 ;
        RECT 2002.330 926.890 2003.510 928.070 ;
        RECT 2002.330 748.490 2003.510 749.670 ;
        RECT 2002.330 746.890 2003.510 748.070 ;
        RECT 2002.330 568.490 2003.510 569.670 ;
        RECT 2002.330 566.890 2003.510 568.070 ;
        RECT 2002.330 388.490 2003.510 389.670 ;
        RECT 2002.330 386.890 2003.510 388.070 ;
        RECT 2002.330 208.490 2003.510 209.670 ;
        RECT 2002.330 206.890 2003.510 208.070 ;
        RECT 2002.330 28.490 2003.510 29.670 ;
        RECT 2002.330 26.890 2003.510 28.070 ;
        RECT 2002.330 -12.110 2003.510 -10.930 ;
        RECT 2002.330 -13.710 2003.510 -12.530 ;
        RECT 2182.330 3532.210 2183.510 3533.390 ;
        RECT 2182.330 3530.610 2183.510 3531.790 ;
        RECT 2182.330 3448.490 2183.510 3449.670 ;
        RECT 2182.330 3446.890 2183.510 3448.070 ;
        RECT 2182.330 3268.490 2183.510 3269.670 ;
        RECT 2182.330 3266.890 2183.510 3268.070 ;
        RECT 2182.330 3088.490 2183.510 3089.670 ;
        RECT 2182.330 3086.890 2183.510 3088.070 ;
        RECT 2182.330 2908.490 2183.510 2909.670 ;
        RECT 2182.330 2906.890 2183.510 2908.070 ;
        RECT 2182.330 2728.490 2183.510 2729.670 ;
        RECT 2182.330 2726.890 2183.510 2728.070 ;
        RECT 2182.330 2548.490 2183.510 2549.670 ;
        RECT 2182.330 2546.890 2183.510 2548.070 ;
        RECT 2182.330 2368.490 2183.510 2369.670 ;
        RECT 2182.330 2366.890 2183.510 2368.070 ;
        RECT 2182.330 2188.490 2183.510 2189.670 ;
        RECT 2182.330 2186.890 2183.510 2188.070 ;
        RECT 2182.330 2008.490 2183.510 2009.670 ;
        RECT 2182.330 2006.890 2183.510 2008.070 ;
        RECT 2182.330 1828.490 2183.510 1829.670 ;
        RECT 2182.330 1826.890 2183.510 1828.070 ;
        RECT 2182.330 1648.490 2183.510 1649.670 ;
        RECT 2182.330 1646.890 2183.510 1648.070 ;
        RECT 2182.330 1468.490 2183.510 1469.670 ;
        RECT 2182.330 1466.890 2183.510 1468.070 ;
        RECT 2182.330 1288.490 2183.510 1289.670 ;
        RECT 2182.330 1286.890 2183.510 1288.070 ;
        RECT 2182.330 1108.490 2183.510 1109.670 ;
        RECT 2182.330 1106.890 2183.510 1108.070 ;
        RECT 2182.330 928.490 2183.510 929.670 ;
        RECT 2182.330 926.890 2183.510 928.070 ;
        RECT 2182.330 748.490 2183.510 749.670 ;
        RECT 2182.330 746.890 2183.510 748.070 ;
        RECT 2182.330 568.490 2183.510 569.670 ;
        RECT 2182.330 566.890 2183.510 568.070 ;
        RECT 2182.330 388.490 2183.510 389.670 ;
        RECT 2182.330 386.890 2183.510 388.070 ;
        RECT 2182.330 208.490 2183.510 209.670 ;
        RECT 2182.330 206.890 2183.510 208.070 ;
        RECT 2182.330 28.490 2183.510 29.670 ;
        RECT 2182.330 26.890 2183.510 28.070 ;
        RECT 2182.330 -12.110 2183.510 -10.930 ;
        RECT 2182.330 -13.710 2183.510 -12.530 ;
        RECT 2362.330 3532.210 2363.510 3533.390 ;
        RECT 2362.330 3530.610 2363.510 3531.790 ;
        RECT 2362.330 3448.490 2363.510 3449.670 ;
        RECT 2362.330 3446.890 2363.510 3448.070 ;
        RECT 2362.330 3268.490 2363.510 3269.670 ;
        RECT 2362.330 3266.890 2363.510 3268.070 ;
        RECT 2362.330 3088.490 2363.510 3089.670 ;
        RECT 2362.330 3086.890 2363.510 3088.070 ;
        RECT 2362.330 2908.490 2363.510 2909.670 ;
        RECT 2362.330 2906.890 2363.510 2908.070 ;
        RECT 2362.330 2728.490 2363.510 2729.670 ;
        RECT 2362.330 2726.890 2363.510 2728.070 ;
        RECT 2362.330 2548.490 2363.510 2549.670 ;
        RECT 2362.330 2546.890 2363.510 2548.070 ;
        RECT 2362.330 2368.490 2363.510 2369.670 ;
        RECT 2362.330 2366.890 2363.510 2368.070 ;
        RECT 2362.330 2188.490 2363.510 2189.670 ;
        RECT 2362.330 2186.890 2363.510 2188.070 ;
        RECT 2362.330 2008.490 2363.510 2009.670 ;
        RECT 2362.330 2006.890 2363.510 2008.070 ;
        RECT 2362.330 1828.490 2363.510 1829.670 ;
        RECT 2362.330 1826.890 2363.510 1828.070 ;
        RECT 2362.330 1648.490 2363.510 1649.670 ;
        RECT 2362.330 1646.890 2363.510 1648.070 ;
        RECT 2362.330 1468.490 2363.510 1469.670 ;
        RECT 2362.330 1466.890 2363.510 1468.070 ;
        RECT 2362.330 1288.490 2363.510 1289.670 ;
        RECT 2362.330 1286.890 2363.510 1288.070 ;
        RECT 2362.330 1108.490 2363.510 1109.670 ;
        RECT 2362.330 1106.890 2363.510 1108.070 ;
        RECT 2362.330 928.490 2363.510 929.670 ;
        RECT 2362.330 926.890 2363.510 928.070 ;
        RECT 2362.330 748.490 2363.510 749.670 ;
        RECT 2362.330 746.890 2363.510 748.070 ;
        RECT 2362.330 568.490 2363.510 569.670 ;
        RECT 2362.330 566.890 2363.510 568.070 ;
        RECT 2362.330 388.490 2363.510 389.670 ;
        RECT 2362.330 386.890 2363.510 388.070 ;
        RECT 2362.330 208.490 2363.510 209.670 ;
        RECT 2362.330 206.890 2363.510 208.070 ;
        RECT 2362.330 28.490 2363.510 29.670 ;
        RECT 2362.330 26.890 2363.510 28.070 ;
        RECT 2362.330 -12.110 2363.510 -10.930 ;
        RECT 2362.330 -13.710 2363.510 -12.530 ;
        RECT 2542.330 3532.210 2543.510 3533.390 ;
        RECT 2542.330 3530.610 2543.510 3531.790 ;
        RECT 2542.330 3448.490 2543.510 3449.670 ;
        RECT 2542.330 3446.890 2543.510 3448.070 ;
        RECT 2542.330 3268.490 2543.510 3269.670 ;
        RECT 2542.330 3266.890 2543.510 3268.070 ;
        RECT 2542.330 3088.490 2543.510 3089.670 ;
        RECT 2542.330 3086.890 2543.510 3088.070 ;
        RECT 2542.330 2908.490 2543.510 2909.670 ;
        RECT 2542.330 2906.890 2543.510 2908.070 ;
        RECT 2542.330 2728.490 2543.510 2729.670 ;
        RECT 2542.330 2726.890 2543.510 2728.070 ;
        RECT 2542.330 2548.490 2543.510 2549.670 ;
        RECT 2542.330 2546.890 2543.510 2548.070 ;
        RECT 2542.330 2368.490 2543.510 2369.670 ;
        RECT 2542.330 2366.890 2543.510 2368.070 ;
        RECT 2542.330 2188.490 2543.510 2189.670 ;
        RECT 2542.330 2186.890 2543.510 2188.070 ;
        RECT 2542.330 2008.490 2543.510 2009.670 ;
        RECT 2542.330 2006.890 2543.510 2008.070 ;
        RECT 2542.330 1828.490 2543.510 1829.670 ;
        RECT 2542.330 1826.890 2543.510 1828.070 ;
        RECT 2542.330 1648.490 2543.510 1649.670 ;
        RECT 2542.330 1646.890 2543.510 1648.070 ;
        RECT 2542.330 1468.490 2543.510 1469.670 ;
        RECT 2542.330 1466.890 2543.510 1468.070 ;
        RECT 2542.330 1288.490 2543.510 1289.670 ;
        RECT 2542.330 1286.890 2543.510 1288.070 ;
        RECT 2542.330 1108.490 2543.510 1109.670 ;
        RECT 2542.330 1106.890 2543.510 1108.070 ;
        RECT 2542.330 928.490 2543.510 929.670 ;
        RECT 2542.330 926.890 2543.510 928.070 ;
        RECT 2542.330 748.490 2543.510 749.670 ;
        RECT 2542.330 746.890 2543.510 748.070 ;
        RECT 2542.330 568.490 2543.510 569.670 ;
        RECT 2542.330 566.890 2543.510 568.070 ;
        RECT 2542.330 388.490 2543.510 389.670 ;
        RECT 2542.330 386.890 2543.510 388.070 ;
        RECT 2542.330 208.490 2543.510 209.670 ;
        RECT 2542.330 206.890 2543.510 208.070 ;
        RECT 2542.330 28.490 2543.510 29.670 ;
        RECT 2542.330 26.890 2543.510 28.070 ;
        RECT 2542.330 -12.110 2543.510 -10.930 ;
        RECT 2542.330 -13.710 2543.510 -12.530 ;
        RECT 2722.330 3532.210 2723.510 3533.390 ;
        RECT 2722.330 3530.610 2723.510 3531.790 ;
        RECT 2722.330 3448.490 2723.510 3449.670 ;
        RECT 2722.330 3446.890 2723.510 3448.070 ;
        RECT 2722.330 3268.490 2723.510 3269.670 ;
        RECT 2722.330 3266.890 2723.510 3268.070 ;
        RECT 2722.330 3088.490 2723.510 3089.670 ;
        RECT 2722.330 3086.890 2723.510 3088.070 ;
        RECT 2722.330 2908.490 2723.510 2909.670 ;
        RECT 2722.330 2906.890 2723.510 2908.070 ;
        RECT 2722.330 2728.490 2723.510 2729.670 ;
        RECT 2722.330 2726.890 2723.510 2728.070 ;
        RECT 2722.330 2548.490 2723.510 2549.670 ;
        RECT 2722.330 2546.890 2723.510 2548.070 ;
        RECT 2722.330 2368.490 2723.510 2369.670 ;
        RECT 2722.330 2366.890 2723.510 2368.070 ;
        RECT 2722.330 2188.490 2723.510 2189.670 ;
        RECT 2722.330 2186.890 2723.510 2188.070 ;
        RECT 2722.330 2008.490 2723.510 2009.670 ;
        RECT 2722.330 2006.890 2723.510 2008.070 ;
        RECT 2722.330 1828.490 2723.510 1829.670 ;
        RECT 2722.330 1826.890 2723.510 1828.070 ;
        RECT 2722.330 1648.490 2723.510 1649.670 ;
        RECT 2722.330 1646.890 2723.510 1648.070 ;
        RECT 2722.330 1468.490 2723.510 1469.670 ;
        RECT 2722.330 1466.890 2723.510 1468.070 ;
        RECT 2722.330 1288.490 2723.510 1289.670 ;
        RECT 2722.330 1286.890 2723.510 1288.070 ;
        RECT 2722.330 1108.490 2723.510 1109.670 ;
        RECT 2722.330 1106.890 2723.510 1108.070 ;
        RECT 2722.330 928.490 2723.510 929.670 ;
        RECT 2722.330 926.890 2723.510 928.070 ;
        RECT 2722.330 748.490 2723.510 749.670 ;
        RECT 2722.330 746.890 2723.510 748.070 ;
        RECT 2722.330 568.490 2723.510 569.670 ;
        RECT 2722.330 566.890 2723.510 568.070 ;
        RECT 2722.330 388.490 2723.510 389.670 ;
        RECT 2722.330 386.890 2723.510 388.070 ;
        RECT 2722.330 208.490 2723.510 209.670 ;
        RECT 2722.330 206.890 2723.510 208.070 ;
        RECT 2722.330 28.490 2723.510 29.670 ;
        RECT 2722.330 26.890 2723.510 28.070 ;
        RECT 2722.330 -12.110 2723.510 -10.930 ;
        RECT 2722.330 -13.710 2723.510 -12.530 ;
        RECT 2902.330 3532.210 2903.510 3533.390 ;
        RECT 2902.330 3530.610 2903.510 3531.790 ;
        RECT 2902.330 3448.490 2903.510 3449.670 ;
        RECT 2902.330 3446.890 2903.510 3448.070 ;
        RECT 2902.330 3268.490 2903.510 3269.670 ;
        RECT 2902.330 3266.890 2903.510 3268.070 ;
        RECT 2902.330 3088.490 2903.510 3089.670 ;
        RECT 2902.330 3086.890 2903.510 3088.070 ;
        RECT 2902.330 2908.490 2903.510 2909.670 ;
        RECT 2902.330 2906.890 2903.510 2908.070 ;
        RECT 2902.330 2728.490 2903.510 2729.670 ;
        RECT 2902.330 2726.890 2903.510 2728.070 ;
        RECT 2902.330 2548.490 2903.510 2549.670 ;
        RECT 2902.330 2546.890 2903.510 2548.070 ;
        RECT 2902.330 2368.490 2903.510 2369.670 ;
        RECT 2902.330 2366.890 2903.510 2368.070 ;
        RECT 2902.330 2188.490 2903.510 2189.670 ;
        RECT 2902.330 2186.890 2903.510 2188.070 ;
        RECT 2902.330 2008.490 2903.510 2009.670 ;
        RECT 2902.330 2006.890 2903.510 2008.070 ;
        RECT 2902.330 1828.490 2903.510 1829.670 ;
        RECT 2902.330 1826.890 2903.510 1828.070 ;
        RECT 2902.330 1648.490 2903.510 1649.670 ;
        RECT 2902.330 1646.890 2903.510 1648.070 ;
        RECT 2902.330 1468.490 2903.510 1469.670 ;
        RECT 2902.330 1466.890 2903.510 1468.070 ;
        RECT 2902.330 1288.490 2903.510 1289.670 ;
        RECT 2902.330 1286.890 2903.510 1288.070 ;
        RECT 2902.330 1108.490 2903.510 1109.670 ;
        RECT 2902.330 1106.890 2903.510 1108.070 ;
        RECT 2902.330 928.490 2903.510 929.670 ;
        RECT 2902.330 926.890 2903.510 928.070 ;
        RECT 2902.330 748.490 2903.510 749.670 ;
        RECT 2902.330 746.890 2903.510 748.070 ;
        RECT 2902.330 568.490 2903.510 569.670 ;
        RECT 2902.330 566.890 2903.510 568.070 ;
        RECT 2902.330 388.490 2903.510 389.670 ;
        RECT 2902.330 386.890 2903.510 388.070 ;
        RECT 2902.330 208.490 2903.510 209.670 ;
        RECT 2902.330 206.890 2903.510 208.070 ;
        RECT 2902.330 28.490 2903.510 29.670 ;
        RECT 2902.330 26.890 2903.510 28.070 ;
        RECT 2902.330 -12.110 2903.510 -10.930 ;
        RECT 2902.330 -13.710 2903.510 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3448.490 2937.890 3449.670 ;
        RECT 2936.710 3446.890 2937.890 3448.070 ;
        RECT 2936.710 3268.490 2937.890 3269.670 ;
        RECT 2936.710 3266.890 2937.890 3268.070 ;
        RECT 2936.710 3088.490 2937.890 3089.670 ;
        RECT 2936.710 3086.890 2937.890 3088.070 ;
        RECT 2936.710 2908.490 2937.890 2909.670 ;
        RECT 2936.710 2906.890 2937.890 2908.070 ;
        RECT 2936.710 2728.490 2937.890 2729.670 ;
        RECT 2936.710 2726.890 2937.890 2728.070 ;
        RECT 2936.710 2548.490 2937.890 2549.670 ;
        RECT 2936.710 2546.890 2937.890 2548.070 ;
        RECT 2936.710 2368.490 2937.890 2369.670 ;
        RECT 2936.710 2366.890 2937.890 2368.070 ;
        RECT 2936.710 2188.490 2937.890 2189.670 ;
        RECT 2936.710 2186.890 2937.890 2188.070 ;
        RECT 2936.710 2008.490 2937.890 2009.670 ;
        RECT 2936.710 2006.890 2937.890 2008.070 ;
        RECT 2936.710 1828.490 2937.890 1829.670 ;
        RECT 2936.710 1826.890 2937.890 1828.070 ;
        RECT 2936.710 1648.490 2937.890 1649.670 ;
        RECT 2936.710 1646.890 2937.890 1648.070 ;
        RECT 2936.710 1468.490 2937.890 1469.670 ;
        RECT 2936.710 1466.890 2937.890 1468.070 ;
        RECT 2936.710 1288.490 2937.890 1289.670 ;
        RECT 2936.710 1286.890 2937.890 1288.070 ;
        RECT 2936.710 1108.490 2937.890 1109.670 ;
        RECT 2936.710 1106.890 2937.890 1108.070 ;
        RECT 2936.710 928.490 2937.890 929.670 ;
        RECT 2936.710 926.890 2937.890 928.070 ;
        RECT 2936.710 748.490 2937.890 749.670 ;
        RECT 2936.710 746.890 2937.890 748.070 ;
        RECT 2936.710 568.490 2937.890 569.670 ;
        RECT 2936.710 566.890 2937.890 568.070 ;
        RECT 2936.710 388.490 2937.890 389.670 ;
        RECT 2936.710 386.890 2937.890 388.070 ;
        RECT 2936.710 208.490 2937.890 209.670 ;
        RECT 2936.710 206.890 2937.890 208.070 ;
        RECT 2936.710 28.490 2937.890 29.670 ;
        RECT 2936.710 26.890 2937.890 28.070 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.130 3533.450 -16.230 3533.510 ;
        RECT 21.470 3533.450 24.370 3533.510 ;
        RECT 201.470 3533.450 204.370 3533.510 ;
        RECT 381.470 3533.450 384.370 3533.510 ;
        RECT 561.470 3533.450 564.370 3533.510 ;
        RECT 741.470 3533.450 744.370 3533.510 ;
        RECT 921.470 3533.450 924.370 3533.510 ;
        RECT 1101.470 3533.450 1104.370 3533.510 ;
        RECT 1281.470 3533.450 1284.370 3533.510 ;
        RECT 1461.470 3533.450 1464.370 3533.510 ;
        RECT 1641.470 3533.450 1644.370 3533.510 ;
        RECT 1821.470 3533.450 1824.370 3533.510 ;
        RECT 2001.470 3533.450 2004.370 3533.510 ;
        RECT 2181.470 3533.450 2184.370 3533.510 ;
        RECT 2361.470 3533.450 2364.370 3533.510 ;
        RECT 2541.470 3533.450 2544.370 3533.510 ;
        RECT 2721.470 3533.450 2724.370 3533.510 ;
        RECT 2901.470 3533.450 2904.370 3533.510 ;
        RECT 2935.850 3533.450 2938.750 3533.510 ;
        RECT -19.130 3530.550 2938.750 3533.450 ;
        RECT -19.130 3530.490 -16.230 3530.550 ;
        RECT 21.470 3530.490 24.370 3530.550 ;
        RECT 201.470 3530.490 204.370 3530.550 ;
        RECT 381.470 3530.490 384.370 3530.550 ;
        RECT 561.470 3530.490 564.370 3530.550 ;
        RECT 741.470 3530.490 744.370 3530.550 ;
        RECT 921.470 3530.490 924.370 3530.550 ;
        RECT 1101.470 3530.490 1104.370 3530.550 ;
        RECT 1281.470 3530.490 1284.370 3530.550 ;
        RECT 1461.470 3530.490 1464.370 3530.550 ;
        RECT 1641.470 3530.490 1644.370 3530.550 ;
        RECT 1821.470 3530.490 1824.370 3530.550 ;
        RECT 2001.470 3530.490 2004.370 3530.550 ;
        RECT 2181.470 3530.490 2184.370 3530.550 ;
        RECT 2361.470 3530.490 2364.370 3530.550 ;
        RECT 2541.470 3530.490 2544.370 3530.550 ;
        RECT 2721.470 3530.490 2724.370 3530.550 ;
        RECT 2901.470 3530.490 2904.370 3530.550 ;
        RECT 2935.850 3530.490 2938.750 3530.550 ;
        RECT -19.130 3449.730 -16.230 3449.790 ;
        RECT 21.470 3449.730 24.370 3449.790 ;
        RECT 201.470 3449.730 204.370 3449.790 ;
        RECT 381.470 3449.730 384.370 3449.790 ;
        RECT 561.470 3449.730 564.370 3449.790 ;
        RECT 741.470 3449.730 744.370 3449.790 ;
        RECT 921.470 3449.730 924.370 3449.790 ;
        RECT 1101.470 3449.730 1104.370 3449.790 ;
        RECT 1281.470 3449.730 1284.370 3449.790 ;
        RECT 1461.470 3449.730 1464.370 3449.790 ;
        RECT 1641.470 3449.730 1644.370 3449.790 ;
        RECT 1821.470 3449.730 1824.370 3449.790 ;
        RECT 2001.470 3449.730 2004.370 3449.790 ;
        RECT 2181.470 3449.730 2184.370 3449.790 ;
        RECT 2361.470 3449.730 2364.370 3449.790 ;
        RECT 2541.470 3449.730 2544.370 3449.790 ;
        RECT 2721.470 3449.730 2724.370 3449.790 ;
        RECT 2901.470 3449.730 2904.370 3449.790 ;
        RECT 2935.850 3449.730 2938.750 3449.790 ;
        RECT -23.730 3446.830 2943.350 3449.730 ;
        RECT -19.130 3446.770 -16.230 3446.830 ;
        RECT 21.470 3446.770 24.370 3446.830 ;
        RECT 201.470 3446.770 204.370 3446.830 ;
        RECT 381.470 3446.770 384.370 3446.830 ;
        RECT 561.470 3446.770 564.370 3446.830 ;
        RECT 741.470 3446.770 744.370 3446.830 ;
        RECT 921.470 3446.770 924.370 3446.830 ;
        RECT 1101.470 3446.770 1104.370 3446.830 ;
        RECT 1281.470 3446.770 1284.370 3446.830 ;
        RECT 1461.470 3446.770 1464.370 3446.830 ;
        RECT 1641.470 3446.770 1644.370 3446.830 ;
        RECT 1821.470 3446.770 1824.370 3446.830 ;
        RECT 2001.470 3446.770 2004.370 3446.830 ;
        RECT 2181.470 3446.770 2184.370 3446.830 ;
        RECT 2361.470 3446.770 2364.370 3446.830 ;
        RECT 2541.470 3446.770 2544.370 3446.830 ;
        RECT 2721.470 3446.770 2724.370 3446.830 ;
        RECT 2901.470 3446.770 2904.370 3446.830 ;
        RECT 2935.850 3446.770 2938.750 3446.830 ;
        RECT -19.130 3269.730 -16.230 3269.790 ;
        RECT 21.470 3269.730 24.370 3269.790 ;
        RECT 201.470 3269.730 204.370 3269.790 ;
        RECT 381.470 3269.730 384.370 3269.790 ;
        RECT 561.470 3269.730 564.370 3269.790 ;
        RECT 741.470 3269.730 744.370 3269.790 ;
        RECT 921.470 3269.730 924.370 3269.790 ;
        RECT 1101.470 3269.730 1104.370 3269.790 ;
        RECT 1281.470 3269.730 1284.370 3269.790 ;
        RECT 1461.470 3269.730 1464.370 3269.790 ;
        RECT 1641.470 3269.730 1644.370 3269.790 ;
        RECT 1821.470 3269.730 1824.370 3269.790 ;
        RECT 2001.470 3269.730 2004.370 3269.790 ;
        RECT 2181.470 3269.730 2184.370 3269.790 ;
        RECT 2361.470 3269.730 2364.370 3269.790 ;
        RECT 2541.470 3269.730 2544.370 3269.790 ;
        RECT 2721.470 3269.730 2724.370 3269.790 ;
        RECT 2901.470 3269.730 2904.370 3269.790 ;
        RECT 2935.850 3269.730 2938.750 3269.790 ;
        RECT -23.730 3266.830 2943.350 3269.730 ;
        RECT -19.130 3266.770 -16.230 3266.830 ;
        RECT 21.470 3266.770 24.370 3266.830 ;
        RECT 201.470 3266.770 204.370 3266.830 ;
        RECT 381.470 3266.770 384.370 3266.830 ;
        RECT 561.470 3266.770 564.370 3266.830 ;
        RECT 741.470 3266.770 744.370 3266.830 ;
        RECT 921.470 3266.770 924.370 3266.830 ;
        RECT 1101.470 3266.770 1104.370 3266.830 ;
        RECT 1281.470 3266.770 1284.370 3266.830 ;
        RECT 1461.470 3266.770 1464.370 3266.830 ;
        RECT 1641.470 3266.770 1644.370 3266.830 ;
        RECT 1821.470 3266.770 1824.370 3266.830 ;
        RECT 2001.470 3266.770 2004.370 3266.830 ;
        RECT 2181.470 3266.770 2184.370 3266.830 ;
        RECT 2361.470 3266.770 2364.370 3266.830 ;
        RECT 2541.470 3266.770 2544.370 3266.830 ;
        RECT 2721.470 3266.770 2724.370 3266.830 ;
        RECT 2901.470 3266.770 2904.370 3266.830 ;
        RECT 2935.850 3266.770 2938.750 3266.830 ;
        RECT -19.130 3089.730 -16.230 3089.790 ;
        RECT 21.470 3089.730 24.370 3089.790 ;
        RECT 201.470 3089.730 204.370 3089.790 ;
        RECT 381.470 3089.730 384.370 3089.790 ;
        RECT 561.470 3089.730 564.370 3089.790 ;
        RECT 741.470 3089.730 744.370 3089.790 ;
        RECT 921.470 3089.730 924.370 3089.790 ;
        RECT 1101.470 3089.730 1104.370 3089.790 ;
        RECT 1281.470 3089.730 1284.370 3089.790 ;
        RECT 1461.470 3089.730 1464.370 3089.790 ;
        RECT 1641.470 3089.730 1644.370 3089.790 ;
        RECT 1821.470 3089.730 1824.370 3089.790 ;
        RECT 2001.470 3089.730 2004.370 3089.790 ;
        RECT 2181.470 3089.730 2184.370 3089.790 ;
        RECT 2361.470 3089.730 2364.370 3089.790 ;
        RECT 2541.470 3089.730 2544.370 3089.790 ;
        RECT 2721.470 3089.730 2724.370 3089.790 ;
        RECT 2901.470 3089.730 2904.370 3089.790 ;
        RECT 2935.850 3089.730 2938.750 3089.790 ;
        RECT -23.730 3086.830 2943.350 3089.730 ;
        RECT -19.130 3086.770 -16.230 3086.830 ;
        RECT 21.470 3086.770 24.370 3086.830 ;
        RECT 201.470 3086.770 204.370 3086.830 ;
        RECT 381.470 3086.770 384.370 3086.830 ;
        RECT 561.470 3086.770 564.370 3086.830 ;
        RECT 741.470 3086.770 744.370 3086.830 ;
        RECT 921.470 3086.770 924.370 3086.830 ;
        RECT 1101.470 3086.770 1104.370 3086.830 ;
        RECT 1281.470 3086.770 1284.370 3086.830 ;
        RECT 1461.470 3086.770 1464.370 3086.830 ;
        RECT 1641.470 3086.770 1644.370 3086.830 ;
        RECT 1821.470 3086.770 1824.370 3086.830 ;
        RECT 2001.470 3086.770 2004.370 3086.830 ;
        RECT 2181.470 3086.770 2184.370 3086.830 ;
        RECT 2361.470 3086.770 2364.370 3086.830 ;
        RECT 2541.470 3086.770 2544.370 3086.830 ;
        RECT 2721.470 3086.770 2724.370 3086.830 ;
        RECT 2901.470 3086.770 2904.370 3086.830 ;
        RECT 2935.850 3086.770 2938.750 3086.830 ;
        RECT -19.130 2909.730 -16.230 2909.790 ;
        RECT 21.470 2909.730 24.370 2909.790 ;
        RECT 201.470 2909.730 204.370 2909.790 ;
        RECT 381.470 2909.730 384.370 2909.790 ;
        RECT 561.470 2909.730 564.370 2909.790 ;
        RECT 741.470 2909.730 744.370 2909.790 ;
        RECT 921.470 2909.730 924.370 2909.790 ;
        RECT 1101.470 2909.730 1104.370 2909.790 ;
        RECT 1281.470 2909.730 1284.370 2909.790 ;
        RECT 1461.470 2909.730 1464.370 2909.790 ;
        RECT 1641.470 2909.730 1644.370 2909.790 ;
        RECT 1821.470 2909.730 1824.370 2909.790 ;
        RECT 2001.470 2909.730 2004.370 2909.790 ;
        RECT 2181.470 2909.730 2184.370 2909.790 ;
        RECT 2361.470 2909.730 2364.370 2909.790 ;
        RECT 2541.470 2909.730 2544.370 2909.790 ;
        RECT 2721.470 2909.730 2724.370 2909.790 ;
        RECT 2901.470 2909.730 2904.370 2909.790 ;
        RECT 2935.850 2909.730 2938.750 2909.790 ;
        RECT -23.730 2906.830 2943.350 2909.730 ;
        RECT -19.130 2906.770 -16.230 2906.830 ;
        RECT 21.470 2906.770 24.370 2906.830 ;
        RECT 201.470 2906.770 204.370 2906.830 ;
        RECT 381.470 2906.770 384.370 2906.830 ;
        RECT 561.470 2906.770 564.370 2906.830 ;
        RECT 741.470 2906.770 744.370 2906.830 ;
        RECT 921.470 2906.770 924.370 2906.830 ;
        RECT 1101.470 2906.770 1104.370 2906.830 ;
        RECT 1281.470 2906.770 1284.370 2906.830 ;
        RECT 1461.470 2906.770 1464.370 2906.830 ;
        RECT 1641.470 2906.770 1644.370 2906.830 ;
        RECT 1821.470 2906.770 1824.370 2906.830 ;
        RECT 2001.470 2906.770 2004.370 2906.830 ;
        RECT 2181.470 2906.770 2184.370 2906.830 ;
        RECT 2361.470 2906.770 2364.370 2906.830 ;
        RECT 2541.470 2906.770 2544.370 2906.830 ;
        RECT 2721.470 2906.770 2724.370 2906.830 ;
        RECT 2901.470 2906.770 2904.370 2906.830 ;
        RECT 2935.850 2906.770 2938.750 2906.830 ;
        RECT -19.130 2729.730 -16.230 2729.790 ;
        RECT 21.470 2729.730 24.370 2729.790 ;
        RECT 201.470 2729.730 204.370 2729.790 ;
        RECT 381.470 2729.730 384.370 2729.790 ;
        RECT 561.470 2729.730 564.370 2729.790 ;
        RECT 741.470 2729.730 744.370 2729.790 ;
        RECT 921.470 2729.730 924.370 2729.790 ;
        RECT 1101.470 2729.730 1104.370 2729.790 ;
        RECT 1281.470 2729.730 1284.370 2729.790 ;
        RECT 1461.470 2729.730 1464.370 2729.790 ;
        RECT 1641.470 2729.730 1644.370 2729.790 ;
        RECT 1821.470 2729.730 1824.370 2729.790 ;
        RECT 2001.470 2729.730 2004.370 2729.790 ;
        RECT 2181.470 2729.730 2184.370 2729.790 ;
        RECT 2361.470 2729.730 2364.370 2729.790 ;
        RECT 2541.470 2729.730 2544.370 2729.790 ;
        RECT 2721.470 2729.730 2724.370 2729.790 ;
        RECT 2901.470 2729.730 2904.370 2729.790 ;
        RECT 2935.850 2729.730 2938.750 2729.790 ;
        RECT -23.730 2726.830 2943.350 2729.730 ;
        RECT -19.130 2726.770 -16.230 2726.830 ;
        RECT 21.470 2726.770 24.370 2726.830 ;
        RECT 201.470 2726.770 204.370 2726.830 ;
        RECT 381.470 2726.770 384.370 2726.830 ;
        RECT 561.470 2726.770 564.370 2726.830 ;
        RECT 741.470 2726.770 744.370 2726.830 ;
        RECT 921.470 2726.770 924.370 2726.830 ;
        RECT 1101.470 2726.770 1104.370 2726.830 ;
        RECT 1281.470 2726.770 1284.370 2726.830 ;
        RECT 1461.470 2726.770 1464.370 2726.830 ;
        RECT 1641.470 2726.770 1644.370 2726.830 ;
        RECT 1821.470 2726.770 1824.370 2726.830 ;
        RECT 2001.470 2726.770 2004.370 2726.830 ;
        RECT 2181.470 2726.770 2184.370 2726.830 ;
        RECT 2361.470 2726.770 2364.370 2726.830 ;
        RECT 2541.470 2726.770 2544.370 2726.830 ;
        RECT 2721.470 2726.770 2724.370 2726.830 ;
        RECT 2901.470 2726.770 2904.370 2726.830 ;
        RECT 2935.850 2726.770 2938.750 2726.830 ;
        RECT -19.130 2549.730 -16.230 2549.790 ;
        RECT 21.470 2549.730 24.370 2549.790 ;
        RECT 201.470 2549.730 204.370 2549.790 ;
        RECT 381.470 2549.730 384.370 2549.790 ;
        RECT 561.470 2549.730 564.370 2549.790 ;
        RECT 741.470 2549.730 744.370 2549.790 ;
        RECT 921.470 2549.730 924.370 2549.790 ;
        RECT 1101.470 2549.730 1104.370 2549.790 ;
        RECT 1281.470 2549.730 1284.370 2549.790 ;
        RECT 1461.470 2549.730 1464.370 2549.790 ;
        RECT 1641.470 2549.730 1644.370 2549.790 ;
        RECT 1821.470 2549.730 1824.370 2549.790 ;
        RECT 2001.470 2549.730 2004.370 2549.790 ;
        RECT 2181.470 2549.730 2184.370 2549.790 ;
        RECT 2361.470 2549.730 2364.370 2549.790 ;
        RECT 2541.470 2549.730 2544.370 2549.790 ;
        RECT 2721.470 2549.730 2724.370 2549.790 ;
        RECT 2901.470 2549.730 2904.370 2549.790 ;
        RECT 2935.850 2549.730 2938.750 2549.790 ;
        RECT -23.730 2546.830 2943.350 2549.730 ;
        RECT -19.130 2546.770 -16.230 2546.830 ;
        RECT 21.470 2546.770 24.370 2546.830 ;
        RECT 201.470 2546.770 204.370 2546.830 ;
        RECT 381.470 2546.770 384.370 2546.830 ;
        RECT 561.470 2546.770 564.370 2546.830 ;
        RECT 741.470 2546.770 744.370 2546.830 ;
        RECT 921.470 2546.770 924.370 2546.830 ;
        RECT 1101.470 2546.770 1104.370 2546.830 ;
        RECT 1281.470 2546.770 1284.370 2546.830 ;
        RECT 1461.470 2546.770 1464.370 2546.830 ;
        RECT 1641.470 2546.770 1644.370 2546.830 ;
        RECT 1821.470 2546.770 1824.370 2546.830 ;
        RECT 2001.470 2546.770 2004.370 2546.830 ;
        RECT 2181.470 2546.770 2184.370 2546.830 ;
        RECT 2361.470 2546.770 2364.370 2546.830 ;
        RECT 2541.470 2546.770 2544.370 2546.830 ;
        RECT 2721.470 2546.770 2724.370 2546.830 ;
        RECT 2901.470 2546.770 2904.370 2546.830 ;
        RECT 2935.850 2546.770 2938.750 2546.830 ;
        RECT -19.130 2369.730 -16.230 2369.790 ;
        RECT 21.470 2369.730 24.370 2369.790 ;
        RECT 201.470 2369.730 204.370 2369.790 ;
        RECT 381.470 2369.730 384.370 2369.790 ;
        RECT 561.470 2369.730 564.370 2369.790 ;
        RECT 741.470 2369.730 744.370 2369.790 ;
        RECT 921.470 2369.730 924.370 2369.790 ;
        RECT 1101.470 2369.730 1104.370 2369.790 ;
        RECT 1281.470 2369.730 1284.370 2369.790 ;
        RECT 1461.470 2369.730 1464.370 2369.790 ;
        RECT 1641.470 2369.730 1644.370 2369.790 ;
        RECT 1821.470 2369.730 1824.370 2369.790 ;
        RECT 2001.470 2369.730 2004.370 2369.790 ;
        RECT 2181.470 2369.730 2184.370 2369.790 ;
        RECT 2361.470 2369.730 2364.370 2369.790 ;
        RECT 2541.470 2369.730 2544.370 2369.790 ;
        RECT 2721.470 2369.730 2724.370 2369.790 ;
        RECT 2901.470 2369.730 2904.370 2369.790 ;
        RECT 2935.850 2369.730 2938.750 2369.790 ;
        RECT -23.730 2366.830 2943.350 2369.730 ;
        RECT -19.130 2366.770 -16.230 2366.830 ;
        RECT 21.470 2366.770 24.370 2366.830 ;
        RECT 201.470 2366.770 204.370 2366.830 ;
        RECT 381.470 2366.770 384.370 2366.830 ;
        RECT 561.470 2366.770 564.370 2366.830 ;
        RECT 741.470 2366.770 744.370 2366.830 ;
        RECT 921.470 2366.770 924.370 2366.830 ;
        RECT 1101.470 2366.770 1104.370 2366.830 ;
        RECT 1281.470 2366.770 1284.370 2366.830 ;
        RECT 1461.470 2366.770 1464.370 2366.830 ;
        RECT 1641.470 2366.770 1644.370 2366.830 ;
        RECT 1821.470 2366.770 1824.370 2366.830 ;
        RECT 2001.470 2366.770 2004.370 2366.830 ;
        RECT 2181.470 2366.770 2184.370 2366.830 ;
        RECT 2361.470 2366.770 2364.370 2366.830 ;
        RECT 2541.470 2366.770 2544.370 2366.830 ;
        RECT 2721.470 2366.770 2724.370 2366.830 ;
        RECT 2901.470 2366.770 2904.370 2366.830 ;
        RECT 2935.850 2366.770 2938.750 2366.830 ;
        RECT -19.130 2189.730 -16.230 2189.790 ;
        RECT 21.470 2189.730 24.370 2189.790 ;
        RECT 201.470 2189.730 204.370 2189.790 ;
        RECT 381.470 2189.730 384.370 2189.790 ;
        RECT 561.470 2189.730 564.370 2189.790 ;
        RECT 741.470 2189.730 744.370 2189.790 ;
        RECT 921.470 2189.730 924.370 2189.790 ;
        RECT 1101.470 2189.730 1104.370 2189.790 ;
        RECT 1281.470 2189.730 1284.370 2189.790 ;
        RECT 1461.470 2189.730 1464.370 2189.790 ;
        RECT 1641.470 2189.730 1644.370 2189.790 ;
        RECT 1821.470 2189.730 1824.370 2189.790 ;
        RECT 2001.470 2189.730 2004.370 2189.790 ;
        RECT 2181.470 2189.730 2184.370 2189.790 ;
        RECT 2361.470 2189.730 2364.370 2189.790 ;
        RECT 2541.470 2189.730 2544.370 2189.790 ;
        RECT 2721.470 2189.730 2724.370 2189.790 ;
        RECT 2901.470 2189.730 2904.370 2189.790 ;
        RECT 2935.850 2189.730 2938.750 2189.790 ;
        RECT -23.730 2186.830 2943.350 2189.730 ;
        RECT -19.130 2186.770 -16.230 2186.830 ;
        RECT 21.470 2186.770 24.370 2186.830 ;
        RECT 201.470 2186.770 204.370 2186.830 ;
        RECT 381.470 2186.770 384.370 2186.830 ;
        RECT 561.470 2186.770 564.370 2186.830 ;
        RECT 741.470 2186.770 744.370 2186.830 ;
        RECT 921.470 2186.770 924.370 2186.830 ;
        RECT 1101.470 2186.770 1104.370 2186.830 ;
        RECT 1281.470 2186.770 1284.370 2186.830 ;
        RECT 1461.470 2186.770 1464.370 2186.830 ;
        RECT 1641.470 2186.770 1644.370 2186.830 ;
        RECT 1821.470 2186.770 1824.370 2186.830 ;
        RECT 2001.470 2186.770 2004.370 2186.830 ;
        RECT 2181.470 2186.770 2184.370 2186.830 ;
        RECT 2361.470 2186.770 2364.370 2186.830 ;
        RECT 2541.470 2186.770 2544.370 2186.830 ;
        RECT 2721.470 2186.770 2724.370 2186.830 ;
        RECT 2901.470 2186.770 2904.370 2186.830 ;
        RECT 2935.850 2186.770 2938.750 2186.830 ;
        RECT -19.130 2009.730 -16.230 2009.790 ;
        RECT 21.470 2009.730 24.370 2009.790 ;
        RECT 201.470 2009.730 204.370 2009.790 ;
        RECT 381.470 2009.730 384.370 2009.790 ;
        RECT 561.470 2009.730 564.370 2009.790 ;
        RECT 741.470 2009.730 744.370 2009.790 ;
        RECT 921.470 2009.730 924.370 2009.790 ;
        RECT 1101.470 2009.730 1104.370 2009.790 ;
        RECT 1281.470 2009.730 1284.370 2009.790 ;
        RECT 1461.470 2009.730 1464.370 2009.790 ;
        RECT 1641.470 2009.730 1644.370 2009.790 ;
        RECT 1821.470 2009.730 1824.370 2009.790 ;
        RECT 2001.470 2009.730 2004.370 2009.790 ;
        RECT 2181.470 2009.730 2184.370 2009.790 ;
        RECT 2361.470 2009.730 2364.370 2009.790 ;
        RECT 2541.470 2009.730 2544.370 2009.790 ;
        RECT 2721.470 2009.730 2724.370 2009.790 ;
        RECT 2901.470 2009.730 2904.370 2009.790 ;
        RECT 2935.850 2009.730 2938.750 2009.790 ;
        RECT -23.730 2006.830 2943.350 2009.730 ;
        RECT -19.130 2006.770 -16.230 2006.830 ;
        RECT 21.470 2006.770 24.370 2006.830 ;
        RECT 201.470 2006.770 204.370 2006.830 ;
        RECT 381.470 2006.770 384.370 2006.830 ;
        RECT 561.470 2006.770 564.370 2006.830 ;
        RECT 741.470 2006.770 744.370 2006.830 ;
        RECT 921.470 2006.770 924.370 2006.830 ;
        RECT 1101.470 2006.770 1104.370 2006.830 ;
        RECT 1281.470 2006.770 1284.370 2006.830 ;
        RECT 1461.470 2006.770 1464.370 2006.830 ;
        RECT 1641.470 2006.770 1644.370 2006.830 ;
        RECT 1821.470 2006.770 1824.370 2006.830 ;
        RECT 2001.470 2006.770 2004.370 2006.830 ;
        RECT 2181.470 2006.770 2184.370 2006.830 ;
        RECT 2361.470 2006.770 2364.370 2006.830 ;
        RECT 2541.470 2006.770 2544.370 2006.830 ;
        RECT 2721.470 2006.770 2724.370 2006.830 ;
        RECT 2901.470 2006.770 2904.370 2006.830 ;
        RECT 2935.850 2006.770 2938.750 2006.830 ;
        RECT -19.130 1829.730 -16.230 1829.790 ;
        RECT 21.470 1829.730 24.370 1829.790 ;
        RECT 201.470 1829.730 204.370 1829.790 ;
        RECT 381.470 1829.730 384.370 1829.790 ;
        RECT 561.470 1829.730 564.370 1829.790 ;
        RECT 741.470 1829.730 744.370 1829.790 ;
        RECT 921.470 1829.730 924.370 1829.790 ;
        RECT 1101.470 1829.730 1104.370 1829.790 ;
        RECT 1281.470 1829.730 1284.370 1829.790 ;
        RECT 1461.470 1829.730 1464.370 1829.790 ;
        RECT 1641.470 1829.730 1644.370 1829.790 ;
        RECT 1821.470 1829.730 1824.370 1829.790 ;
        RECT 2001.470 1829.730 2004.370 1829.790 ;
        RECT 2181.470 1829.730 2184.370 1829.790 ;
        RECT 2361.470 1829.730 2364.370 1829.790 ;
        RECT 2541.470 1829.730 2544.370 1829.790 ;
        RECT 2721.470 1829.730 2724.370 1829.790 ;
        RECT 2901.470 1829.730 2904.370 1829.790 ;
        RECT 2935.850 1829.730 2938.750 1829.790 ;
        RECT -23.730 1826.830 2943.350 1829.730 ;
        RECT -19.130 1826.770 -16.230 1826.830 ;
        RECT 21.470 1826.770 24.370 1826.830 ;
        RECT 201.470 1826.770 204.370 1826.830 ;
        RECT 381.470 1826.770 384.370 1826.830 ;
        RECT 561.470 1826.770 564.370 1826.830 ;
        RECT 741.470 1826.770 744.370 1826.830 ;
        RECT 921.470 1826.770 924.370 1826.830 ;
        RECT 1101.470 1826.770 1104.370 1826.830 ;
        RECT 1281.470 1826.770 1284.370 1826.830 ;
        RECT 1461.470 1826.770 1464.370 1826.830 ;
        RECT 1641.470 1826.770 1644.370 1826.830 ;
        RECT 1821.470 1826.770 1824.370 1826.830 ;
        RECT 2001.470 1826.770 2004.370 1826.830 ;
        RECT 2181.470 1826.770 2184.370 1826.830 ;
        RECT 2361.470 1826.770 2364.370 1826.830 ;
        RECT 2541.470 1826.770 2544.370 1826.830 ;
        RECT 2721.470 1826.770 2724.370 1826.830 ;
        RECT 2901.470 1826.770 2904.370 1826.830 ;
        RECT 2935.850 1826.770 2938.750 1826.830 ;
        RECT -19.130 1649.730 -16.230 1649.790 ;
        RECT 21.470 1649.730 24.370 1649.790 ;
        RECT 201.470 1649.730 204.370 1649.790 ;
        RECT 381.470 1649.730 384.370 1649.790 ;
        RECT 561.470 1649.730 564.370 1649.790 ;
        RECT 741.470 1649.730 744.370 1649.790 ;
        RECT 921.470 1649.730 924.370 1649.790 ;
        RECT 1101.470 1649.730 1104.370 1649.790 ;
        RECT 1281.470 1649.730 1284.370 1649.790 ;
        RECT 1461.470 1649.730 1464.370 1649.790 ;
        RECT 1641.470 1649.730 1644.370 1649.790 ;
        RECT 1821.470 1649.730 1824.370 1649.790 ;
        RECT 2001.470 1649.730 2004.370 1649.790 ;
        RECT 2181.470 1649.730 2184.370 1649.790 ;
        RECT 2361.470 1649.730 2364.370 1649.790 ;
        RECT 2541.470 1649.730 2544.370 1649.790 ;
        RECT 2721.470 1649.730 2724.370 1649.790 ;
        RECT 2901.470 1649.730 2904.370 1649.790 ;
        RECT 2935.850 1649.730 2938.750 1649.790 ;
        RECT -23.730 1646.830 2943.350 1649.730 ;
        RECT -19.130 1646.770 -16.230 1646.830 ;
        RECT 21.470 1646.770 24.370 1646.830 ;
        RECT 201.470 1646.770 204.370 1646.830 ;
        RECT 381.470 1646.770 384.370 1646.830 ;
        RECT 561.470 1646.770 564.370 1646.830 ;
        RECT 741.470 1646.770 744.370 1646.830 ;
        RECT 921.470 1646.770 924.370 1646.830 ;
        RECT 1101.470 1646.770 1104.370 1646.830 ;
        RECT 1281.470 1646.770 1284.370 1646.830 ;
        RECT 1461.470 1646.770 1464.370 1646.830 ;
        RECT 1641.470 1646.770 1644.370 1646.830 ;
        RECT 1821.470 1646.770 1824.370 1646.830 ;
        RECT 2001.470 1646.770 2004.370 1646.830 ;
        RECT 2181.470 1646.770 2184.370 1646.830 ;
        RECT 2361.470 1646.770 2364.370 1646.830 ;
        RECT 2541.470 1646.770 2544.370 1646.830 ;
        RECT 2721.470 1646.770 2724.370 1646.830 ;
        RECT 2901.470 1646.770 2904.370 1646.830 ;
        RECT 2935.850 1646.770 2938.750 1646.830 ;
        RECT -19.130 1469.730 -16.230 1469.790 ;
        RECT 21.470 1469.730 24.370 1469.790 ;
        RECT 201.470 1469.730 204.370 1469.790 ;
        RECT 381.470 1469.730 384.370 1469.790 ;
        RECT 561.470 1469.730 564.370 1469.790 ;
        RECT 741.470 1469.730 744.370 1469.790 ;
        RECT 921.470 1469.730 924.370 1469.790 ;
        RECT 1101.470 1469.730 1104.370 1469.790 ;
        RECT 1281.470 1469.730 1284.370 1469.790 ;
        RECT 1461.470 1469.730 1464.370 1469.790 ;
        RECT 1641.470 1469.730 1644.370 1469.790 ;
        RECT 1821.470 1469.730 1824.370 1469.790 ;
        RECT 2001.470 1469.730 2004.370 1469.790 ;
        RECT 2181.470 1469.730 2184.370 1469.790 ;
        RECT 2361.470 1469.730 2364.370 1469.790 ;
        RECT 2541.470 1469.730 2544.370 1469.790 ;
        RECT 2721.470 1469.730 2724.370 1469.790 ;
        RECT 2901.470 1469.730 2904.370 1469.790 ;
        RECT 2935.850 1469.730 2938.750 1469.790 ;
        RECT -23.730 1466.830 2943.350 1469.730 ;
        RECT -19.130 1466.770 -16.230 1466.830 ;
        RECT 21.470 1466.770 24.370 1466.830 ;
        RECT 201.470 1466.770 204.370 1466.830 ;
        RECT 381.470 1466.770 384.370 1466.830 ;
        RECT 561.470 1466.770 564.370 1466.830 ;
        RECT 741.470 1466.770 744.370 1466.830 ;
        RECT 921.470 1466.770 924.370 1466.830 ;
        RECT 1101.470 1466.770 1104.370 1466.830 ;
        RECT 1281.470 1466.770 1284.370 1466.830 ;
        RECT 1461.470 1466.770 1464.370 1466.830 ;
        RECT 1641.470 1466.770 1644.370 1466.830 ;
        RECT 1821.470 1466.770 1824.370 1466.830 ;
        RECT 2001.470 1466.770 2004.370 1466.830 ;
        RECT 2181.470 1466.770 2184.370 1466.830 ;
        RECT 2361.470 1466.770 2364.370 1466.830 ;
        RECT 2541.470 1466.770 2544.370 1466.830 ;
        RECT 2721.470 1466.770 2724.370 1466.830 ;
        RECT 2901.470 1466.770 2904.370 1466.830 ;
        RECT 2935.850 1466.770 2938.750 1466.830 ;
        RECT -19.130 1289.730 -16.230 1289.790 ;
        RECT 21.470 1289.730 24.370 1289.790 ;
        RECT 201.470 1289.730 204.370 1289.790 ;
        RECT 381.470 1289.730 384.370 1289.790 ;
        RECT 561.470 1289.730 564.370 1289.790 ;
        RECT 741.470 1289.730 744.370 1289.790 ;
        RECT 921.470 1289.730 924.370 1289.790 ;
        RECT 1101.470 1289.730 1104.370 1289.790 ;
        RECT 1281.470 1289.730 1284.370 1289.790 ;
        RECT 1461.470 1289.730 1464.370 1289.790 ;
        RECT 1641.470 1289.730 1644.370 1289.790 ;
        RECT 1821.470 1289.730 1824.370 1289.790 ;
        RECT 2001.470 1289.730 2004.370 1289.790 ;
        RECT 2181.470 1289.730 2184.370 1289.790 ;
        RECT 2361.470 1289.730 2364.370 1289.790 ;
        RECT 2541.470 1289.730 2544.370 1289.790 ;
        RECT 2721.470 1289.730 2724.370 1289.790 ;
        RECT 2901.470 1289.730 2904.370 1289.790 ;
        RECT 2935.850 1289.730 2938.750 1289.790 ;
        RECT -23.730 1286.830 2943.350 1289.730 ;
        RECT -19.130 1286.770 -16.230 1286.830 ;
        RECT 21.470 1286.770 24.370 1286.830 ;
        RECT 201.470 1286.770 204.370 1286.830 ;
        RECT 381.470 1286.770 384.370 1286.830 ;
        RECT 561.470 1286.770 564.370 1286.830 ;
        RECT 741.470 1286.770 744.370 1286.830 ;
        RECT 921.470 1286.770 924.370 1286.830 ;
        RECT 1101.470 1286.770 1104.370 1286.830 ;
        RECT 1281.470 1286.770 1284.370 1286.830 ;
        RECT 1461.470 1286.770 1464.370 1286.830 ;
        RECT 1641.470 1286.770 1644.370 1286.830 ;
        RECT 1821.470 1286.770 1824.370 1286.830 ;
        RECT 2001.470 1286.770 2004.370 1286.830 ;
        RECT 2181.470 1286.770 2184.370 1286.830 ;
        RECT 2361.470 1286.770 2364.370 1286.830 ;
        RECT 2541.470 1286.770 2544.370 1286.830 ;
        RECT 2721.470 1286.770 2724.370 1286.830 ;
        RECT 2901.470 1286.770 2904.370 1286.830 ;
        RECT 2935.850 1286.770 2938.750 1286.830 ;
        RECT -19.130 1109.730 -16.230 1109.790 ;
        RECT 21.470 1109.730 24.370 1109.790 ;
        RECT 201.470 1109.730 204.370 1109.790 ;
        RECT 381.470 1109.730 384.370 1109.790 ;
        RECT 561.470 1109.730 564.370 1109.790 ;
        RECT 741.470 1109.730 744.370 1109.790 ;
        RECT 921.470 1109.730 924.370 1109.790 ;
        RECT 1101.470 1109.730 1104.370 1109.790 ;
        RECT 1281.470 1109.730 1284.370 1109.790 ;
        RECT 1461.470 1109.730 1464.370 1109.790 ;
        RECT 1641.470 1109.730 1644.370 1109.790 ;
        RECT 1821.470 1109.730 1824.370 1109.790 ;
        RECT 2001.470 1109.730 2004.370 1109.790 ;
        RECT 2181.470 1109.730 2184.370 1109.790 ;
        RECT 2361.470 1109.730 2364.370 1109.790 ;
        RECT 2541.470 1109.730 2544.370 1109.790 ;
        RECT 2721.470 1109.730 2724.370 1109.790 ;
        RECT 2901.470 1109.730 2904.370 1109.790 ;
        RECT 2935.850 1109.730 2938.750 1109.790 ;
        RECT -23.730 1106.830 2943.350 1109.730 ;
        RECT -19.130 1106.770 -16.230 1106.830 ;
        RECT 21.470 1106.770 24.370 1106.830 ;
        RECT 201.470 1106.770 204.370 1106.830 ;
        RECT 381.470 1106.770 384.370 1106.830 ;
        RECT 561.470 1106.770 564.370 1106.830 ;
        RECT 741.470 1106.770 744.370 1106.830 ;
        RECT 921.470 1106.770 924.370 1106.830 ;
        RECT 1101.470 1106.770 1104.370 1106.830 ;
        RECT 1281.470 1106.770 1284.370 1106.830 ;
        RECT 1461.470 1106.770 1464.370 1106.830 ;
        RECT 1641.470 1106.770 1644.370 1106.830 ;
        RECT 1821.470 1106.770 1824.370 1106.830 ;
        RECT 2001.470 1106.770 2004.370 1106.830 ;
        RECT 2181.470 1106.770 2184.370 1106.830 ;
        RECT 2361.470 1106.770 2364.370 1106.830 ;
        RECT 2541.470 1106.770 2544.370 1106.830 ;
        RECT 2721.470 1106.770 2724.370 1106.830 ;
        RECT 2901.470 1106.770 2904.370 1106.830 ;
        RECT 2935.850 1106.770 2938.750 1106.830 ;
        RECT -19.130 929.730 -16.230 929.790 ;
        RECT 21.470 929.730 24.370 929.790 ;
        RECT 201.470 929.730 204.370 929.790 ;
        RECT 381.470 929.730 384.370 929.790 ;
        RECT 561.470 929.730 564.370 929.790 ;
        RECT 741.470 929.730 744.370 929.790 ;
        RECT 921.470 929.730 924.370 929.790 ;
        RECT 1101.470 929.730 1104.370 929.790 ;
        RECT 1281.470 929.730 1284.370 929.790 ;
        RECT 1461.470 929.730 1464.370 929.790 ;
        RECT 1641.470 929.730 1644.370 929.790 ;
        RECT 1821.470 929.730 1824.370 929.790 ;
        RECT 2001.470 929.730 2004.370 929.790 ;
        RECT 2181.470 929.730 2184.370 929.790 ;
        RECT 2361.470 929.730 2364.370 929.790 ;
        RECT 2541.470 929.730 2544.370 929.790 ;
        RECT 2721.470 929.730 2724.370 929.790 ;
        RECT 2901.470 929.730 2904.370 929.790 ;
        RECT 2935.850 929.730 2938.750 929.790 ;
        RECT -23.730 926.830 2943.350 929.730 ;
        RECT -19.130 926.770 -16.230 926.830 ;
        RECT 21.470 926.770 24.370 926.830 ;
        RECT 201.470 926.770 204.370 926.830 ;
        RECT 381.470 926.770 384.370 926.830 ;
        RECT 561.470 926.770 564.370 926.830 ;
        RECT 741.470 926.770 744.370 926.830 ;
        RECT 921.470 926.770 924.370 926.830 ;
        RECT 1101.470 926.770 1104.370 926.830 ;
        RECT 1281.470 926.770 1284.370 926.830 ;
        RECT 1461.470 926.770 1464.370 926.830 ;
        RECT 1641.470 926.770 1644.370 926.830 ;
        RECT 1821.470 926.770 1824.370 926.830 ;
        RECT 2001.470 926.770 2004.370 926.830 ;
        RECT 2181.470 926.770 2184.370 926.830 ;
        RECT 2361.470 926.770 2364.370 926.830 ;
        RECT 2541.470 926.770 2544.370 926.830 ;
        RECT 2721.470 926.770 2724.370 926.830 ;
        RECT 2901.470 926.770 2904.370 926.830 ;
        RECT 2935.850 926.770 2938.750 926.830 ;
        RECT -19.130 749.730 -16.230 749.790 ;
        RECT 21.470 749.730 24.370 749.790 ;
        RECT 201.470 749.730 204.370 749.790 ;
        RECT 381.470 749.730 384.370 749.790 ;
        RECT 561.470 749.730 564.370 749.790 ;
        RECT 741.470 749.730 744.370 749.790 ;
        RECT 921.470 749.730 924.370 749.790 ;
        RECT 1101.470 749.730 1104.370 749.790 ;
        RECT 1281.470 749.730 1284.370 749.790 ;
        RECT 1461.470 749.730 1464.370 749.790 ;
        RECT 1641.470 749.730 1644.370 749.790 ;
        RECT 1821.470 749.730 1824.370 749.790 ;
        RECT 2001.470 749.730 2004.370 749.790 ;
        RECT 2181.470 749.730 2184.370 749.790 ;
        RECT 2361.470 749.730 2364.370 749.790 ;
        RECT 2541.470 749.730 2544.370 749.790 ;
        RECT 2721.470 749.730 2724.370 749.790 ;
        RECT 2901.470 749.730 2904.370 749.790 ;
        RECT 2935.850 749.730 2938.750 749.790 ;
        RECT -23.730 746.830 2943.350 749.730 ;
        RECT -19.130 746.770 -16.230 746.830 ;
        RECT 21.470 746.770 24.370 746.830 ;
        RECT 201.470 746.770 204.370 746.830 ;
        RECT 381.470 746.770 384.370 746.830 ;
        RECT 561.470 746.770 564.370 746.830 ;
        RECT 741.470 746.770 744.370 746.830 ;
        RECT 921.470 746.770 924.370 746.830 ;
        RECT 1101.470 746.770 1104.370 746.830 ;
        RECT 1281.470 746.770 1284.370 746.830 ;
        RECT 1461.470 746.770 1464.370 746.830 ;
        RECT 1641.470 746.770 1644.370 746.830 ;
        RECT 1821.470 746.770 1824.370 746.830 ;
        RECT 2001.470 746.770 2004.370 746.830 ;
        RECT 2181.470 746.770 2184.370 746.830 ;
        RECT 2361.470 746.770 2364.370 746.830 ;
        RECT 2541.470 746.770 2544.370 746.830 ;
        RECT 2721.470 746.770 2724.370 746.830 ;
        RECT 2901.470 746.770 2904.370 746.830 ;
        RECT 2935.850 746.770 2938.750 746.830 ;
        RECT -19.130 569.730 -16.230 569.790 ;
        RECT 21.470 569.730 24.370 569.790 ;
        RECT 201.470 569.730 204.370 569.790 ;
        RECT 381.470 569.730 384.370 569.790 ;
        RECT 561.470 569.730 564.370 569.790 ;
        RECT 741.470 569.730 744.370 569.790 ;
        RECT 921.470 569.730 924.370 569.790 ;
        RECT 1101.470 569.730 1104.370 569.790 ;
        RECT 1281.470 569.730 1284.370 569.790 ;
        RECT 1461.470 569.730 1464.370 569.790 ;
        RECT 1641.470 569.730 1644.370 569.790 ;
        RECT 1821.470 569.730 1824.370 569.790 ;
        RECT 2001.470 569.730 2004.370 569.790 ;
        RECT 2181.470 569.730 2184.370 569.790 ;
        RECT 2361.470 569.730 2364.370 569.790 ;
        RECT 2541.470 569.730 2544.370 569.790 ;
        RECT 2721.470 569.730 2724.370 569.790 ;
        RECT 2901.470 569.730 2904.370 569.790 ;
        RECT 2935.850 569.730 2938.750 569.790 ;
        RECT -23.730 566.830 2943.350 569.730 ;
        RECT -19.130 566.770 -16.230 566.830 ;
        RECT 21.470 566.770 24.370 566.830 ;
        RECT 201.470 566.770 204.370 566.830 ;
        RECT 381.470 566.770 384.370 566.830 ;
        RECT 561.470 566.770 564.370 566.830 ;
        RECT 741.470 566.770 744.370 566.830 ;
        RECT 921.470 566.770 924.370 566.830 ;
        RECT 1101.470 566.770 1104.370 566.830 ;
        RECT 1281.470 566.770 1284.370 566.830 ;
        RECT 1461.470 566.770 1464.370 566.830 ;
        RECT 1641.470 566.770 1644.370 566.830 ;
        RECT 1821.470 566.770 1824.370 566.830 ;
        RECT 2001.470 566.770 2004.370 566.830 ;
        RECT 2181.470 566.770 2184.370 566.830 ;
        RECT 2361.470 566.770 2364.370 566.830 ;
        RECT 2541.470 566.770 2544.370 566.830 ;
        RECT 2721.470 566.770 2724.370 566.830 ;
        RECT 2901.470 566.770 2904.370 566.830 ;
        RECT 2935.850 566.770 2938.750 566.830 ;
        RECT -19.130 389.730 -16.230 389.790 ;
        RECT 21.470 389.730 24.370 389.790 ;
        RECT 201.470 389.730 204.370 389.790 ;
        RECT 381.470 389.730 384.370 389.790 ;
        RECT 561.470 389.730 564.370 389.790 ;
        RECT 741.470 389.730 744.370 389.790 ;
        RECT 921.470 389.730 924.370 389.790 ;
        RECT 1101.470 389.730 1104.370 389.790 ;
        RECT 1281.470 389.730 1284.370 389.790 ;
        RECT 1461.470 389.730 1464.370 389.790 ;
        RECT 1641.470 389.730 1644.370 389.790 ;
        RECT 1821.470 389.730 1824.370 389.790 ;
        RECT 2001.470 389.730 2004.370 389.790 ;
        RECT 2181.470 389.730 2184.370 389.790 ;
        RECT 2361.470 389.730 2364.370 389.790 ;
        RECT 2541.470 389.730 2544.370 389.790 ;
        RECT 2721.470 389.730 2724.370 389.790 ;
        RECT 2901.470 389.730 2904.370 389.790 ;
        RECT 2935.850 389.730 2938.750 389.790 ;
        RECT -23.730 386.830 2943.350 389.730 ;
        RECT -19.130 386.770 -16.230 386.830 ;
        RECT 21.470 386.770 24.370 386.830 ;
        RECT 201.470 386.770 204.370 386.830 ;
        RECT 381.470 386.770 384.370 386.830 ;
        RECT 561.470 386.770 564.370 386.830 ;
        RECT 741.470 386.770 744.370 386.830 ;
        RECT 921.470 386.770 924.370 386.830 ;
        RECT 1101.470 386.770 1104.370 386.830 ;
        RECT 1281.470 386.770 1284.370 386.830 ;
        RECT 1461.470 386.770 1464.370 386.830 ;
        RECT 1641.470 386.770 1644.370 386.830 ;
        RECT 1821.470 386.770 1824.370 386.830 ;
        RECT 2001.470 386.770 2004.370 386.830 ;
        RECT 2181.470 386.770 2184.370 386.830 ;
        RECT 2361.470 386.770 2364.370 386.830 ;
        RECT 2541.470 386.770 2544.370 386.830 ;
        RECT 2721.470 386.770 2724.370 386.830 ;
        RECT 2901.470 386.770 2904.370 386.830 ;
        RECT 2935.850 386.770 2938.750 386.830 ;
        RECT -19.130 209.730 -16.230 209.790 ;
        RECT 21.470 209.730 24.370 209.790 ;
        RECT 201.470 209.730 204.370 209.790 ;
        RECT 381.470 209.730 384.370 209.790 ;
        RECT 561.470 209.730 564.370 209.790 ;
        RECT 741.470 209.730 744.370 209.790 ;
        RECT 921.470 209.730 924.370 209.790 ;
        RECT 1101.470 209.730 1104.370 209.790 ;
        RECT 1281.470 209.730 1284.370 209.790 ;
        RECT 1461.470 209.730 1464.370 209.790 ;
        RECT 1641.470 209.730 1644.370 209.790 ;
        RECT 1821.470 209.730 1824.370 209.790 ;
        RECT 2001.470 209.730 2004.370 209.790 ;
        RECT 2181.470 209.730 2184.370 209.790 ;
        RECT 2361.470 209.730 2364.370 209.790 ;
        RECT 2541.470 209.730 2544.370 209.790 ;
        RECT 2721.470 209.730 2724.370 209.790 ;
        RECT 2901.470 209.730 2904.370 209.790 ;
        RECT 2935.850 209.730 2938.750 209.790 ;
        RECT -23.730 206.830 2943.350 209.730 ;
        RECT -19.130 206.770 -16.230 206.830 ;
        RECT 21.470 206.770 24.370 206.830 ;
        RECT 201.470 206.770 204.370 206.830 ;
        RECT 381.470 206.770 384.370 206.830 ;
        RECT 561.470 206.770 564.370 206.830 ;
        RECT 741.470 206.770 744.370 206.830 ;
        RECT 921.470 206.770 924.370 206.830 ;
        RECT 1101.470 206.770 1104.370 206.830 ;
        RECT 1281.470 206.770 1284.370 206.830 ;
        RECT 1461.470 206.770 1464.370 206.830 ;
        RECT 1641.470 206.770 1644.370 206.830 ;
        RECT 1821.470 206.770 1824.370 206.830 ;
        RECT 2001.470 206.770 2004.370 206.830 ;
        RECT 2181.470 206.770 2184.370 206.830 ;
        RECT 2361.470 206.770 2364.370 206.830 ;
        RECT 2541.470 206.770 2544.370 206.830 ;
        RECT 2721.470 206.770 2724.370 206.830 ;
        RECT 2901.470 206.770 2904.370 206.830 ;
        RECT 2935.850 206.770 2938.750 206.830 ;
        RECT -19.130 29.730 -16.230 29.790 ;
        RECT 21.470 29.730 24.370 29.790 ;
        RECT 201.470 29.730 204.370 29.790 ;
        RECT 381.470 29.730 384.370 29.790 ;
        RECT 561.470 29.730 564.370 29.790 ;
        RECT 741.470 29.730 744.370 29.790 ;
        RECT 921.470 29.730 924.370 29.790 ;
        RECT 1101.470 29.730 1104.370 29.790 ;
        RECT 1281.470 29.730 1284.370 29.790 ;
        RECT 1461.470 29.730 1464.370 29.790 ;
        RECT 1641.470 29.730 1644.370 29.790 ;
        RECT 1821.470 29.730 1824.370 29.790 ;
        RECT 2001.470 29.730 2004.370 29.790 ;
        RECT 2181.470 29.730 2184.370 29.790 ;
        RECT 2361.470 29.730 2364.370 29.790 ;
        RECT 2541.470 29.730 2544.370 29.790 ;
        RECT 2721.470 29.730 2724.370 29.790 ;
        RECT 2901.470 29.730 2904.370 29.790 ;
        RECT 2935.850 29.730 2938.750 29.790 ;
        RECT -23.730 26.830 2943.350 29.730 ;
        RECT -19.130 26.770 -16.230 26.830 ;
        RECT 21.470 26.770 24.370 26.830 ;
        RECT 201.470 26.770 204.370 26.830 ;
        RECT 381.470 26.770 384.370 26.830 ;
        RECT 561.470 26.770 564.370 26.830 ;
        RECT 741.470 26.770 744.370 26.830 ;
        RECT 921.470 26.770 924.370 26.830 ;
        RECT 1101.470 26.770 1104.370 26.830 ;
        RECT 1281.470 26.770 1284.370 26.830 ;
        RECT 1461.470 26.770 1464.370 26.830 ;
        RECT 1641.470 26.770 1644.370 26.830 ;
        RECT 1821.470 26.770 1824.370 26.830 ;
        RECT 2001.470 26.770 2004.370 26.830 ;
        RECT 2181.470 26.770 2184.370 26.830 ;
        RECT 2361.470 26.770 2364.370 26.830 ;
        RECT 2541.470 26.770 2544.370 26.830 ;
        RECT 2721.470 26.770 2724.370 26.830 ;
        RECT 2901.470 26.770 2904.370 26.830 ;
        RECT 2935.850 26.770 2938.750 26.830 ;
        RECT -19.130 -10.870 -16.230 -10.810 ;
        RECT 21.470 -10.870 24.370 -10.810 ;
        RECT 201.470 -10.870 204.370 -10.810 ;
        RECT 381.470 -10.870 384.370 -10.810 ;
        RECT 561.470 -10.870 564.370 -10.810 ;
        RECT 741.470 -10.870 744.370 -10.810 ;
        RECT 921.470 -10.870 924.370 -10.810 ;
        RECT 1101.470 -10.870 1104.370 -10.810 ;
        RECT 1281.470 -10.870 1284.370 -10.810 ;
        RECT 1461.470 -10.870 1464.370 -10.810 ;
        RECT 1641.470 -10.870 1644.370 -10.810 ;
        RECT 1821.470 -10.870 1824.370 -10.810 ;
        RECT 2001.470 -10.870 2004.370 -10.810 ;
        RECT 2181.470 -10.870 2184.370 -10.810 ;
        RECT 2361.470 -10.870 2364.370 -10.810 ;
        RECT 2541.470 -10.870 2544.370 -10.810 ;
        RECT 2721.470 -10.870 2724.370 -10.810 ;
        RECT 2901.470 -10.870 2904.370 -10.810 ;
        RECT 2935.850 -10.870 2938.750 -10.810 ;
        RECT -19.130 -13.770 2938.750 -10.870 ;
        RECT -19.130 -13.830 -16.230 -13.770 ;
        RECT 21.470 -13.830 24.370 -13.770 ;
        RECT 201.470 -13.830 204.370 -13.770 ;
        RECT 381.470 -13.830 384.370 -13.770 ;
        RECT 561.470 -13.830 564.370 -13.770 ;
        RECT 741.470 -13.830 744.370 -13.770 ;
        RECT 921.470 -13.830 924.370 -13.770 ;
        RECT 1101.470 -13.830 1104.370 -13.770 ;
        RECT 1281.470 -13.830 1284.370 -13.770 ;
        RECT 1461.470 -13.830 1464.370 -13.770 ;
        RECT 1641.470 -13.830 1644.370 -13.770 ;
        RECT 1821.470 -13.830 1824.370 -13.770 ;
        RECT 2001.470 -13.830 2004.370 -13.770 ;
        RECT 2181.470 -13.830 2184.370 -13.770 ;
        RECT 2361.470 -13.830 2364.370 -13.770 ;
        RECT 2541.470 -13.830 2544.370 -13.770 ;
        RECT 2721.470 -13.830 2724.370 -13.770 ;
        RECT 2901.470 -13.830 2904.370 -13.770 ;
        RECT 2935.850 -13.830 2938.750 -13.770 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.730 -18.370 -20.830 3538.050 ;
        RECT 111.470 -18.370 114.370 3538.050 ;
        RECT 291.470 -18.370 294.370 3538.050 ;
        RECT 471.470 -18.370 474.370 3538.050 ;
        RECT 651.470 -18.370 654.370 3538.050 ;
        RECT 831.470 -18.370 834.370 3538.050 ;
        RECT 1011.470 -18.370 1014.370 3538.050 ;
        RECT 1191.470 -18.370 1194.370 3538.050 ;
        RECT 1371.470 -18.370 1374.370 3538.050 ;
        RECT 1551.470 -18.370 1554.370 3538.050 ;
        RECT 1731.470 -18.370 1734.370 3538.050 ;
        RECT 1911.470 -18.370 1914.370 3538.050 ;
        RECT 2091.470 -18.370 2094.370 3538.050 ;
        RECT 2271.470 -18.370 2274.370 3538.050 ;
        RECT 2451.470 -18.370 2454.370 3538.050 ;
        RECT 2631.470 -18.370 2634.370 3538.050 ;
        RECT 2811.470 -18.370 2814.370 3538.050 ;
        RECT 2940.450 -18.370 2943.350 3538.050 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3358.490 -21.690 3359.670 ;
        RECT -22.870 3356.890 -21.690 3358.070 ;
        RECT -22.870 3178.490 -21.690 3179.670 ;
        RECT -22.870 3176.890 -21.690 3178.070 ;
        RECT -22.870 2998.490 -21.690 2999.670 ;
        RECT -22.870 2996.890 -21.690 2998.070 ;
        RECT -22.870 2818.490 -21.690 2819.670 ;
        RECT -22.870 2816.890 -21.690 2818.070 ;
        RECT -22.870 2638.490 -21.690 2639.670 ;
        RECT -22.870 2636.890 -21.690 2638.070 ;
        RECT -22.870 2458.490 -21.690 2459.670 ;
        RECT -22.870 2456.890 -21.690 2458.070 ;
        RECT -22.870 2278.490 -21.690 2279.670 ;
        RECT -22.870 2276.890 -21.690 2278.070 ;
        RECT -22.870 2098.490 -21.690 2099.670 ;
        RECT -22.870 2096.890 -21.690 2098.070 ;
        RECT -22.870 1918.490 -21.690 1919.670 ;
        RECT -22.870 1916.890 -21.690 1918.070 ;
        RECT -22.870 1738.490 -21.690 1739.670 ;
        RECT -22.870 1736.890 -21.690 1738.070 ;
        RECT -22.870 1558.490 -21.690 1559.670 ;
        RECT -22.870 1556.890 -21.690 1558.070 ;
        RECT -22.870 1378.490 -21.690 1379.670 ;
        RECT -22.870 1376.890 -21.690 1378.070 ;
        RECT -22.870 1198.490 -21.690 1199.670 ;
        RECT -22.870 1196.890 -21.690 1198.070 ;
        RECT -22.870 1018.490 -21.690 1019.670 ;
        RECT -22.870 1016.890 -21.690 1018.070 ;
        RECT -22.870 838.490 -21.690 839.670 ;
        RECT -22.870 836.890 -21.690 838.070 ;
        RECT -22.870 658.490 -21.690 659.670 ;
        RECT -22.870 656.890 -21.690 658.070 ;
        RECT -22.870 478.490 -21.690 479.670 ;
        RECT -22.870 476.890 -21.690 478.070 ;
        RECT -22.870 298.490 -21.690 299.670 ;
        RECT -22.870 296.890 -21.690 298.070 ;
        RECT -22.870 118.490 -21.690 119.670 ;
        RECT -22.870 116.890 -21.690 118.070 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.330 3536.810 113.510 3537.990 ;
        RECT 112.330 3535.210 113.510 3536.390 ;
        RECT 112.330 3358.490 113.510 3359.670 ;
        RECT 112.330 3356.890 113.510 3358.070 ;
        RECT 112.330 3178.490 113.510 3179.670 ;
        RECT 112.330 3176.890 113.510 3178.070 ;
        RECT 112.330 2998.490 113.510 2999.670 ;
        RECT 112.330 2996.890 113.510 2998.070 ;
        RECT 112.330 2818.490 113.510 2819.670 ;
        RECT 112.330 2816.890 113.510 2818.070 ;
        RECT 112.330 2638.490 113.510 2639.670 ;
        RECT 112.330 2636.890 113.510 2638.070 ;
        RECT 112.330 2458.490 113.510 2459.670 ;
        RECT 112.330 2456.890 113.510 2458.070 ;
        RECT 112.330 2278.490 113.510 2279.670 ;
        RECT 112.330 2276.890 113.510 2278.070 ;
        RECT 112.330 2098.490 113.510 2099.670 ;
        RECT 112.330 2096.890 113.510 2098.070 ;
        RECT 112.330 1918.490 113.510 1919.670 ;
        RECT 112.330 1916.890 113.510 1918.070 ;
        RECT 112.330 1738.490 113.510 1739.670 ;
        RECT 112.330 1736.890 113.510 1738.070 ;
        RECT 112.330 1558.490 113.510 1559.670 ;
        RECT 112.330 1556.890 113.510 1558.070 ;
        RECT 112.330 1378.490 113.510 1379.670 ;
        RECT 112.330 1376.890 113.510 1378.070 ;
        RECT 112.330 1198.490 113.510 1199.670 ;
        RECT 112.330 1196.890 113.510 1198.070 ;
        RECT 112.330 1018.490 113.510 1019.670 ;
        RECT 112.330 1016.890 113.510 1018.070 ;
        RECT 112.330 838.490 113.510 839.670 ;
        RECT 112.330 836.890 113.510 838.070 ;
        RECT 112.330 658.490 113.510 659.670 ;
        RECT 112.330 656.890 113.510 658.070 ;
        RECT 112.330 478.490 113.510 479.670 ;
        RECT 112.330 476.890 113.510 478.070 ;
        RECT 112.330 298.490 113.510 299.670 ;
        RECT 112.330 296.890 113.510 298.070 ;
        RECT 112.330 118.490 113.510 119.670 ;
        RECT 112.330 116.890 113.510 118.070 ;
        RECT 112.330 -16.710 113.510 -15.530 ;
        RECT 112.330 -18.310 113.510 -17.130 ;
        RECT 292.330 3536.810 293.510 3537.990 ;
        RECT 292.330 3535.210 293.510 3536.390 ;
        RECT 292.330 3358.490 293.510 3359.670 ;
        RECT 292.330 3356.890 293.510 3358.070 ;
        RECT 292.330 3178.490 293.510 3179.670 ;
        RECT 292.330 3176.890 293.510 3178.070 ;
        RECT 292.330 2998.490 293.510 2999.670 ;
        RECT 292.330 2996.890 293.510 2998.070 ;
        RECT 292.330 2818.490 293.510 2819.670 ;
        RECT 292.330 2816.890 293.510 2818.070 ;
        RECT 292.330 2638.490 293.510 2639.670 ;
        RECT 292.330 2636.890 293.510 2638.070 ;
        RECT 292.330 2458.490 293.510 2459.670 ;
        RECT 292.330 2456.890 293.510 2458.070 ;
        RECT 292.330 2278.490 293.510 2279.670 ;
        RECT 292.330 2276.890 293.510 2278.070 ;
        RECT 292.330 2098.490 293.510 2099.670 ;
        RECT 292.330 2096.890 293.510 2098.070 ;
        RECT 292.330 1918.490 293.510 1919.670 ;
        RECT 292.330 1916.890 293.510 1918.070 ;
        RECT 292.330 1738.490 293.510 1739.670 ;
        RECT 292.330 1736.890 293.510 1738.070 ;
        RECT 292.330 1558.490 293.510 1559.670 ;
        RECT 292.330 1556.890 293.510 1558.070 ;
        RECT 292.330 1378.490 293.510 1379.670 ;
        RECT 292.330 1376.890 293.510 1378.070 ;
        RECT 292.330 1198.490 293.510 1199.670 ;
        RECT 292.330 1196.890 293.510 1198.070 ;
        RECT 292.330 1018.490 293.510 1019.670 ;
        RECT 292.330 1016.890 293.510 1018.070 ;
        RECT 292.330 838.490 293.510 839.670 ;
        RECT 292.330 836.890 293.510 838.070 ;
        RECT 292.330 658.490 293.510 659.670 ;
        RECT 292.330 656.890 293.510 658.070 ;
        RECT 292.330 478.490 293.510 479.670 ;
        RECT 292.330 476.890 293.510 478.070 ;
        RECT 292.330 298.490 293.510 299.670 ;
        RECT 292.330 296.890 293.510 298.070 ;
        RECT 292.330 118.490 293.510 119.670 ;
        RECT 292.330 116.890 293.510 118.070 ;
        RECT 292.330 -16.710 293.510 -15.530 ;
        RECT 292.330 -18.310 293.510 -17.130 ;
        RECT 472.330 3536.810 473.510 3537.990 ;
        RECT 472.330 3535.210 473.510 3536.390 ;
        RECT 472.330 3358.490 473.510 3359.670 ;
        RECT 472.330 3356.890 473.510 3358.070 ;
        RECT 472.330 3178.490 473.510 3179.670 ;
        RECT 472.330 3176.890 473.510 3178.070 ;
        RECT 472.330 2998.490 473.510 2999.670 ;
        RECT 472.330 2996.890 473.510 2998.070 ;
        RECT 472.330 2818.490 473.510 2819.670 ;
        RECT 472.330 2816.890 473.510 2818.070 ;
        RECT 472.330 2638.490 473.510 2639.670 ;
        RECT 472.330 2636.890 473.510 2638.070 ;
        RECT 472.330 2458.490 473.510 2459.670 ;
        RECT 472.330 2456.890 473.510 2458.070 ;
        RECT 472.330 2278.490 473.510 2279.670 ;
        RECT 472.330 2276.890 473.510 2278.070 ;
        RECT 472.330 2098.490 473.510 2099.670 ;
        RECT 472.330 2096.890 473.510 2098.070 ;
        RECT 472.330 1918.490 473.510 1919.670 ;
        RECT 472.330 1916.890 473.510 1918.070 ;
        RECT 472.330 1738.490 473.510 1739.670 ;
        RECT 472.330 1736.890 473.510 1738.070 ;
        RECT 472.330 1558.490 473.510 1559.670 ;
        RECT 472.330 1556.890 473.510 1558.070 ;
        RECT 472.330 1378.490 473.510 1379.670 ;
        RECT 472.330 1376.890 473.510 1378.070 ;
        RECT 472.330 1198.490 473.510 1199.670 ;
        RECT 472.330 1196.890 473.510 1198.070 ;
        RECT 472.330 1018.490 473.510 1019.670 ;
        RECT 472.330 1016.890 473.510 1018.070 ;
        RECT 472.330 838.490 473.510 839.670 ;
        RECT 472.330 836.890 473.510 838.070 ;
        RECT 472.330 658.490 473.510 659.670 ;
        RECT 472.330 656.890 473.510 658.070 ;
        RECT 472.330 478.490 473.510 479.670 ;
        RECT 472.330 476.890 473.510 478.070 ;
        RECT 472.330 298.490 473.510 299.670 ;
        RECT 472.330 296.890 473.510 298.070 ;
        RECT 472.330 118.490 473.510 119.670 ;
        RECT 472.330 116.890 473.510 118.070 ;
        RECT 472.330 -16.710 473.510 -15.530 ;
        RECT 472.330 -18.310 473.510 -17.130 ;
        RECT 652.330 3536.810 653.510 3537.990 ;
        RECT 652.330 3535.210 653.510 3536.390 ;
        RECT 652.330 3358.490 653.510 3359.670 ;
        RECT 652.330 3356.890 653.510 3358.070 ;
        RECT 652.330 3178.490 653.510 3179.670 ;
        RECT 652.330 3176.890 653.510 3178.070 ;
        RECT 652.330 2998.490 653.510 2999.670 ;
        RECT 652.330 2996.890 653.510 2998.070 ;
        RECT 652.330 2818.490 653.510 2819.670 ;
        RECT 652.330 2816.890 653.510 2818.070 ;
        RECT 652.330 2638.490 653.510 2639.670 ;
        RECT 652.330 2636.890 653.510 2638.070 ;
        RECT 652.330 2458.490 653.510 2459.670 ;
        RECT 652.330 2456.890 653.510 2458.070 ;
        RECT 652.330 2278.490 653.510 2279.670 ;
        RECT 652.330 2276.890 653.510 2278.070 ;
        RECT 652.330 2098.490 653.510 2099.670 ;
        RECT 652.330 2096.890 653.510 2098.070 ;
        RECT 652.330 1918.490 653.510 1919.670 ;
        RECT 652.330 1916.890 653.510 1918.070 ;
        RECT 652.330 1738.490 653.510 1739.670 ;
        RECT 652.330 1736.890 653.510 1738.070 ;
        RECT 652.330 1558.490 653.510 1559.670 ;
        RECT 652.330 1556.890 653.510 1558.070 ;
        RECT 652.330 1378.490 653.510 1379.670 ;
        RECT 652.330 1376.890 653.510 1378.070 ;
        RECT 652.330 1198.490 653.510 1199.670 ;
        RECT 652.330 1196.890 653.510 1198.070 ;
        RECT 652.330 1018.490 653.510 1019.670 ;
        RECT 652.330 1016.890 653.510 1018.070 ;
        RECT 652.330 838.490 653.510 839.670 ;
        RECT 652.330 836.890 653.510 838.070 ;
        RECT 652.330 658.490 653.510 659.670 ;
        RECT 652.330 656.890 653.510 658.070 ;
        RECT 652.330 478.490 653.510 479.670 ;
        RECT 652.330 476.890 653.510 478.070 ;
        RECT 652.330 298.490 653.510 299.670 ;
        RECT 652.330 296.890 653.510 298.070 ;
        RECT 652.330 118.490 653.510 119.670 ;
        RECT 652.330 116.890 653.510 118.070 ;
        RECT 652.330 -16.710 653.510 -15.530 ;
        RECT 652.330 -18.310 653.510 -17.130 ;
        RECT 832.330 3536.810 833.510 3537.990 ;
        RECT 832.330 3535.210 833.510 3536.390 ;
        RECT 832.330 3358.490 833.510 3359.670 ;
        RECT 832.330 3356.890 833.510 3358.070 ;
        RECT 832.330 3178.490 833.510 3179.670 ;
        RECT 832.330 3176.890 833.510 3178.070 ;
        RECT 832.330 2998.490 833.510 2999.670 ;
        RECT 832.330 2996.890 833.510 2998.070 ;
        RECT 832.330 2818.490 833.510 2819.670 ;
        RECT 832.330 2816.890 833.510 2818.070 ;
        RECT 832.330 2638.490 833.510 2639.670 ;
        RECT 832.330 2636.890 833.510 2638.070 ;
        RECT 832.330 2458.490 833.510 2459.670 ;
        RECT 832.330 2456.890 833.510 2458.070 ;
        RECT 832.330 2278.490 833.510 2279.670 ;
        RECT 832.330 2276.890 833.510 2278.070 ;
        RECT 832.330 2098.490 833.510 2099.670 ;
        RECT 832.330 2096.890 833.510 2098.070 ;
        RECT 832.330 1918.490 833.510 1919.670 ;
        RECT 832.330 1916.890 833.510 1918.070 ;
        RECT 832.330 1738.490 833.510 1739.670 ;
        RECT 832.330 1736.890 833.510 1738.070 ;
        RECT 832.330 1558.490 833.510 1559.670 ;
        RECT 832.330 1556.890 833.510 1558.070 ;
        RECT 832.330 1378.490 833.510 1379.670 ;
        RECT 832.330 1376.890 833.510 1378.070 ;
        RECT 832.330 1198.490 833.510 1199.670 ;
        RECT 832.330 1196.890 833.510 1198.070 ;
        RECT 832.330 1018.490 833.510 1019.670 ;
        RECT 832.330 1016.890 833.510 1018.070 ;
        RECT 832.330 838.490 833.510 839.670 ;
        RECT 832.330 836.890 833.510 838.070 ;
        RECT 832.330 658.490 833.510 659.670 ;
        RECT 832.330 656.890 833.510 658.070 ;
        RECT 832.330 478.490 833.510 479.670 ;
        RECT 832.330 476.890 833.510 478.070 ;
        RECT 832.330 298.490 833.510 299.670 ;
        RECT 832.330 296.890 833.510 298.070 ;
        RECT 832.330 118.490 833.510 119.670 ;
        RECT 832.330 116.890 833.510 118.070 ;
        RECT 832.330 -16.710 833.510 -15.530 ;
        RECT 832.330 -18.310 833.510 -17.130 ;
        RECT 1012.330 3536.810 1013.510 3537.990 ;
        RECT 1012.330 3535.210 1013.510 3536.390 ;
        RECT 1012.330 3358.490 1013.510 3359.670 ;
        RECT 1012.330 3356.890 1013.510 3358.070 ;
        RECT 1012.330 3178.490 1013.510 3179.670 ;
        RECT 1012.330 3176.890 1013.510 3178.070 ;
        RECT 1012.330 2998.490 1013.510 2999.670 ;
        RECT 1012.330 2996.890 1013.510 2998.070 ;
        RECT 1012.330 2818.490 1013.510 2819.670 ;
        RECT 1012.330 2816.890 1013.510 2818.070 ;
        RECT 1012.330 2638.490 1013.510 2639.670 ;
        RECT 1012.330 2636.890 1013.510 2638.070 ;
        RECT 1012.330 2458.490 1013.510 2459.670 ;
        RECT 1012.330 2456.890 1013.510 2458.070 ;
        RECT 1012.330 2278.490 1013.510 2279.670 ;
        RECT 1012.330 2276.890 1013.510 2278.070 ;
        RECT 1012.330 2098.490 1013.510 2099.670 ;
        RECT 1012.330 2096.890 1013.510 2098.070 ;
        RECT 1012.330 1918.490 1013.510 1919.670 ;
        RECT 1012.330 1916.890 1013.510 1918.070 ;
        RECT 1012.330 1738.490 1013.510 1739.670 ;
        RECT 1012.330 1736.890 1013.510 1738.070 ;
        RECT 1012.330 1558.490 1013.510 1559.670 ;
        RECT 1012.330 1556.890 1013.510 1558.070 ;
        RECT 1012.330 1378.490 1013.510 1379.670 ;
        RECT 1012.330 1376.890 1013.510 1378.070 ;
        RECT 1012.330 1198.490 1013.510 1199.670 ;
        RECT 1012.330 1196.890 1013.510 1198.070 ;
        RECT 1012.330 1018.490 1013.510 1019.670 ;
        RECT 1012.330 1016.890 1013.510 1018.070 ;
        RECT 1012.330 838.490 1013.510 839.670 ;
        RECT 1012.330 836.890 1013.510 838.070 ;
        RECT 1012.330 658.490 1013.510 659.670 ;
        RECT 1012.330 656.890 1013.510 658.070 ;
        RECT 1012.330 478.490 1013.510 479.670 ;
        RECT 1012.330 476.890 1013.510 478.070 ;
        RECT 1012.330 298.490 1013.510 299.670 ;
        RECT 1012.330 296.890 1013.510 298.070 ;
        RECT 1012.330 118.490 1013.510 119.670 ;
        RECT 1012.330 116.890 1013.510 118.070 ;
        RECT 1012.330 -16.710 1013.510 -15.530 ;
        RECT 1012.330 -18.310 1013.510 -17.130 ;
        RECT 1192.330 3536.810 1193.510 3537.990 ;
        RECT 1192.330 3535.210 1193.510 3536.390 ;
        RECT 1192.330 3358.490 1193.510 3359.670 ;
        RECT 1192.330 3356.890 1193.510 3358.070 ;
        RECT 1192.330 3178.490 1193.510 3179.670 ;
        RECT 1192.330 3176.890 1193.510 3178.070 ;
        RECT 1192.330 2998.490 1193.510 2999.670 ;
        RECT 1192.330 2996.890 1193.510 2998.070 ;
        RECT 1192.330 2818.490 1193.510 2819.670 ;
        RECT 1192.330 2816.890 1193.510 2818.070 ;
        RECT 1192.330 2638.490 1193.510 2639.670 ;
        RECT 1192.330 2636.890 1193.510 2638.070 ;
        RECT 1192.330 2458.490 1193.510 2459.670 ;
        RECT 1192.330 2456.890 1193.510 2458.070 ;
        RECT 1192.330 2278.490 1193.510 2279.670 ;
        RECT 1192.330 2276.890 1193.510 2278.070 ;
        RECT 1192.330 2098.490 1193.510 2099.670 ;
        RECT 1192.330 2096.890 1193.510 2098.070 ;
        RECT 1192.330 1918.490 1193.510 1919.670 ;
        RECT 1192.330 1916.890 1193.510 1918.070 ;
        RECT 1192.330 1738.490 1193.510 1739.670 ;
        RECT 1192.330 1736.890 1193.510 1738.070 ;
        RECT 1192.330 1558.490 1193.510 1559.670 ;
        RECT 1192.330 1556.890 1193.510 1558.070 ;
        RECT 1192.330 1378.490 1193.510 1379.670 ;
        RECT 1192.330 1376.890 1193.510 1378.070 ;
        RECT 1192.330 1198.490 1193.510 1199.670 ;
        RECT 1192.330 1196.890 1193.510 1198.070 ;
        RECT 1192.330 1018.490 1193.510 1019.670 ;
        RECT 1192.330 1016.890 1193.510 1018.070 ;
        RECT 1192.330 838.490 1193.510 839.670 ;
        RECT 1192.330 836.890 1193.510 838.070 ;
        RECT 1192.330 658.490 1193.510 659.670 ;
        RECT 1192.330 656.890 1193.510 658.070 ;
        RECT 1192.330 478.490 1193.510 479.670 ;
        RECT 1192.330 476.890 1193.510 478.070 ;
        RECT 1192.330 298.490 1193.510 299.670 ;
        RECT 1192.330 296.890 1193.510 298.070 ;
        RECT 1192.330 118.490 1193.510 119.670 ;
        RECT 1192.330 116.890 1193.510 118.070 ;
        RECT 1192.330 -16.710 1193.510 -15.530 ;
        RECT 1192.330 -18.310 1193.510 -17.130 ;
        RECT 1372.330 3536.810 1373.510 3537.990 ;
        RECT 1372.330 3535.210 1373.510 3536.390 ;
        RECT 1372.330 3358.490 1373.510 3359.670 ;
        RECT 1372.330 3356.890 1373.510 3358.070 ;
        RECT 1372.330 3178.490 1373.510 3179.670 ;
        RECT 1372.330 3176.890 1373.510 3178.070 ;
        RECT 1372.330 2998.490 1373.510 2999.670 ;
        RECT 1372.330 2996.890 1373.510 2998.070 ;
        RECT 1372.330 2818.490 1373.510 2819.670 ;
        RECT 1372.330 2816.890 1373.510 2818.070 ;
        RECT 1372.330 2638.490 1373.510 2639.670 ;
        RECT 1372.330 2636.890 1373.510 2638.070 ;
        RECT 1372.330 2458.490 1373.510 2459.670 ;
        RECT 1372.330 2456.890 1373.510 2458.070 ;
        RECT 1372.330 2278.490 1373.510 2279.670 ;
        RECT 1372.330 2276.890 1373.510 2278.070 ;
        RECT 1372.330 2098.490 1373.510 2099.670 ;
        RECT 1372.330 2096.890 1373.510 2098.070 ;
        RECT 1372.330 1918.490 1373.510 1919.670 ;
        RECT 1372.330 1916.890 1373.510 1918.070 ;
        RECT 1372.330 1738.490 1373.510 1739.670 ;
        RECT 1372.330 1736.890 1373.510 1738.070 ;
        RECT 1372.330 1558.490 1373.510 1559.670 ;
        RECT 1372.330 1556.890 1373.510 1558.070 ;
        RECT 1372.330 1378.490 1373.510 1379.670 ;
        RECT 1372.330 1376.890 1373.510 1378.070 ;
        RECT 1372.330 1198.490 1373.510 1199.670 ;
        RECT 1372.330 1196.890 1373.510 1198.070 ;
        RECT 1372.330 1018.490 1373.510 1019.670 ;
        RECT 1372.330 1016.890 1373.510 1018.070 ;
        RECT 1372.330 838.490 1373.510 839.670 ;
        RECT 1372.330 836.890 1373.510 838.070 ;
        RECT 1372.330 658.490 1373.510 659.670 ;
        RECT 1372.330 656.890 1373.510 658.070 ;
        RECT 1372.330 478.490 1373.510 479.670 ;
        RECT 1372.330 476.890 1373.510 478.070 ;
        RECT 1372.330 298.490 1373.510 299.670 ;
        RECT 1372.330 296.890 1373.510 298.070 ;
        RECT 1372.330 118.490 1373.510 119.670 ;
        RECT 1372.330 116.890 1373.510 118.070 ;
        RECT 1372.330 -16.710 1373.510 -15.530 ;
        RECT 1372.330 -18.310 1373.510 -17.130 ;
        RECT 1552.330 3536.810 1553.510 3537.990 ;
        RECT 1552.330 3535.210 1553.510 3536.390 ;
        RECT 1552.330 3358.490 1553.510 3359.670 ;
        RECT 1552.330 3356.890 1553.510 3358.070 ;
        RECT 1552.330 3178.490 1553.510 3179.670 ;
        RECT 1552.330 3176.890 1553.510 3178.070 ;
        RECT 1552.330 2998.490 1553.510 2999.670 ;
        RECT 1552.330 2996.890 1553.510 2998.070 ;
        RECT 1552.330 2818.490 1553.510 2819.670 ;
        RECT 1552.330 2816.890 1553.510 2818.070 ;
        RECT 1552.330 2638.490 1553.510 2639.670 ;
        RECT 1552.330 2636.890 1553.510 2638.070 ;
        RECT 1552.330 2458.490 1553.510 2459.670 ;
        RECT 1552.330 2456.890 1553.510 2458.070 ;
        RECT 1552.330 2278.490 1553.510 2279.670 ;
        RECT 1552.330 2276.890 1553.510 2278.070 ;
        RECT 1552.330 2098.490 1553.510 2099.670 ;
        RECT 1552.330 2096.890 1553.510 2098.070 ;
        RECT 1552.330 1918.490 1553.510 1919.670 ;
        RECT 1552.330 1916.890 1553.510 1918.070 ;
        RECT 1552.330 1738.490 1553.510 1739.670 ;
        RECT 1552.330 1736.890 1553.510 1738.070 ;
        RECT 1552.330 1558.490 1553.510 1559.670 ;
        RECT 1552.330 1556.890 1553.510 1558.070 ;
        RECT 1552.330 1378.490 1553.510 1379.670 ;
        RECT 1552.330 1376.890 1553.510 1378.070 ;
        RECT 1552.330 1198.490 1553.510 1199.670 ;
        RECT 1552.330 1196.890 1553.510 1198.070 ;
        RECT 1552.330 1018.490 1553.510 1019.670 ;
        RECT 1552.330 1016.890 1553.510 1018.070 ;
        RECT 1552.330 838.490 1553.510 839.670 ;
        RECT 1552.330 836.890 1553.510 838.070 ;
        RECT 1552.330 658.490 1553.510 659.670 ;
        RECT 1552.330 656.890 1553.510 658.070 ;
        RECT 1552.330 478.490 1553.510 479.670 ;
        RECT 1552.330 476.890 1553.510 478.070 ;
        RECT 1552.330 298.490 1553.510 299.670 ;
        RECT 1552.330 296.890 1553.510 298.070 ;
        RECT 1552.330 118.490 1553.510 119.670 ;
        RECT 1552.330 116.890 1553.510 118.070 ;
        RECT 1552.330 -16.710 1553.510 -15.530 ;
        RECT 1552.330 -18.310 1553.510 -17.130 ;
        RECT 1732.330 3536.810 1733.510 3537.990 ;
        RECT 1732.330 3535.210 1733.510 3536.390 ;
        RECT 1732.330 3358.490 1733.510 3359.670 ;
        RECT 1732.330 3356.890 1733.510 3358.070 ;
        RECT 1732.330 3178.490 1733.510 3179.670 ;
        RECT 1732.330 3176.890 1733.510 3178.070 ;
        RECT 1732.330 2998.490 1733.510 2999.670 ;
        RECT 1732.330 2996.890 1733.510 2998.070 ;
        RECT 1732.330 2818.490 1733.510 2819.670 ;
        RECT 1732.330 2816.890 1733.510 2818.070 ;
        RECT 1732.330 2638.490 1733.510 2639.670 ;
        RECT 1732.330 2636.890 1733.510 2638.070 ;
        RECT 1732.330 2458.490 1733.510 2459.670 ;
        RECT 1732.330 2456.890 1733.510 2458.070 ;
        RECT 1732.330 2278.490 1733.510 2279.670 ;
        RECT 1732.330 2276.890 1733.510 2278.070 ;
        RECT 1732.330 2098.490 1733.510 2099.670 ;
        RECT 1732.330 2096.890 1733.510 2098.070 ;
        RECT 1732.330 1918.490 1733.510 1919.670 ;
        RECT 1732.330 1916.890 1733.510 1918.070 ;
        RECT 1732.330 1738.490 1733.510 1739.670 ;
        RECT 1732.330 1736.890 1733.510 1738.070 ;
        RECT 1732.330 1558.490 1733.510 1559.670 ;
        RECT 1732.330 1556.890 1733.510 1558.070 ;
        RECT 1732.330 1378.490 1733.510 1379.670 ;
        RECT 1732.330 1376.890 1733.510 1378.070 ;
        RECT 1732.330 1198.490 1733.510 1199.670 ;
        RECT 1732.330 1196.890 1733.510 1198.070 ;
        RECT 1732.330 1018.490 1733.510 1019.670 ;
        RECT 1732.330 1016.890 1733.510 1018.070 ;
        RECT 1732.330 838.490 1733.510 839.670 ;
        RECT 1732.330 836.890 1733.510 838.070 ;
        RECT 1732.330 658.490 1733.510 659.670 ;
        RECT 1732.330 656.890 1733.510 658.070 ;
        RECT 1732.330 478.490 1733.510 479.670 ;
        RECT 1732.330 476.890 1733.510 478.070 ;
        RECT 1732.330 298.490 1733.510 299.670 ;
        RECT 1732.330 296.890 1733.510 298.070 ;
        RECT 1732.330 118.490 1733.510 119.670 ;
        RECT 1732.330 116.890 1733.510 118.070 ;
        RECT 1732.330 -16.710 1733.510 -15.530 ;
        RECT 1732.330 -18.310 1733.510 -17.130 ;
        RECT 1912.330 3536.810 1913.510 3537.990 ;
        RECT 1912.330 3535.210 1913.510 3536.390 ;
        RECT 1912.330 3358.490 1913.510 3359.670 ;
        RECT 1912.330 3356.890 1913.510 3358.070 ;
        RECT 1912.330 3178.490 1913.510 3179.670 ;
        RECT 1912.330 3176.890 1913.510 3178.070 ;
        RECT 1912.330 2998.490 1913.510 2999.670 ;
        RECT 1912.330 2996.890 1913.510 2998.070 ;
        RECT 1912.330 2818.490 1913.510 2819.670 ;
        RECT 1912.330 2816.890 1913.510 2818.070 ;
        RECT 1912.330 2638.490 1913.510 2639.670 ;
        RECT 1912.330 2636.890 1913.510 2638.070 ;
        RECT 1912.330 2458.490 1913.510 2459.670 ;
        RECT 1912.330 2456.890 1913.510 2458.070 ;
        RECT 1912.330 2278.490 1913.510 2279.670 ;
        RECT 1912.330 2276.890 1913.510 2278.070 ;
        RECT 1912.330 2098.490 1913.510 2099.670 ;
        RECT 1912.330 2096.890 1913.510 2098.070 ;
        RECT 1912.330 1918.490 1913.510 1919.670 ;
        RECT 1912.330 1916.890 1913.510 1918.070 ;
        RECT 1912.330 1738.490 1913.510 1739.670 ;
        RECT 1912.330 1736.890 1913.510 1738.070 ;
        RECT 1912.330 1558.490 1913.510 1559.670 ;
        RECT 1912.330 1556.890 1913.510 1558.070 ;
        RECT 1912.330 1378.490 1913.510 1379.670 ;
        RECT 1912.330 1376.890 1913.510 1378.070 ;
        RECT 1912.330 1198.490 1913.510 1199.670 ;
        RECT 1912.330 1196.890 1913.510 1198.070 ;
        RECT 1912.330 1018.490 1913.510 1019.670 ;
        RECT 1912.330 1016.890 1913.510 1018.070 ;
        RECT 1912.330 838.490 1913.510 839.670 ;
        RECT 1912.330 836.890 1913.510 838.070 ;
        RECT 1912.330 658.490 1913.510 659.670 ;
        RECT 1912.330 656.890 1913.510 658.070 ;
        RECT 1912.330 478.490 1913.510 479.670 ;
        RECT 1912.330 476.890 1913.510 478.070 ;
        RECT 1912.330 298.490 1913.510 299.670 ;
        RECT 1912.330 296.890 1913.510 298.070 ;
        RECT 1912.330 118.490 1913.510 119.670 ;
        RECT 1912.330 116.890 1913.510 118.070 ;
        RECT 1912.330 -16.710 1913.510 -15.530 ;
        RECT 1912.330 -18.310 1913.510 -17.130 ;
        RECT 2092.330 3536.810 2093.510 3537.990 ;
        RECT 2092.330 3535.210 2093.510 3536.390 ;
        RECT 2092.330 3358.490 2093.510 3359.670 ;
        RECT 2092.330 3356.890 2093.510 3358.070 ;
        RECT 2092.330 3178.490 2093.510 3179.670 ;
        RECT 2092.330 3176.890 2093.510 3178.070 ;
        RECT 2092.330 2998.490 2093.510 2999.670 ;
        RECT 2092.330 2996.890 2093.510 2998.070 ;
        RECT 2092.330 2818.490 2093.510 2819.670 ;
        RECT 2092.330 2816.890 2093.510 2818.070 ;
        RECT 2092.330 2638.490 2093.510 2639.670 ;
        RECT 2092.330 2636.890 2093.510 2638.070 ;
        RECT 2092.330 2458.490 2093.510 2459.670 ;
        RECT 2092.330 2456.890 2093.510 2458.070 ;
        RECT 2092.330 2278.490 2093.510 2279.670 ;
        RECT 2092.330 2276.890 2093.510 2278.070 ;
        RECT 2092.330 2098.490 2093.510 2099.670 ;
        RECT 2092.330 2096.890 2093.510 2098.070 ;
        RECT 2092.330 1918.490 2093.510 1919.670 ;
        RECT 2092.330 1916.890 2093.510 1918.070 ;
        RECT 2092.330 1738.490 2093.510 1739.670 ;
        RECT 2092.330 1736.890 2093.510 1738.070 ;
        RECT 2092.330 1558.490 2093.510 1559.670 ;
        RECT 2092.330 1556.890 2093.510 1558.070 ;
        RECT 2092.330 1378.490 2093.510 1379.670 ;
        RECT 2092.330 1376.890 2093.510 1378.070 ;
        RECT 2092.330 1198.490 2093.510 1199.670 ;
        RECT 2092.330 1196.890 2093.510 1198.070 ;
        RECT 2092.330 1018.490 2093.510 1019.670 ;
        RECT 2092.330 1016.890 2093.510 1018.070 ;
        RECT 2092.330 838.490 2093.510 839.670 ;
        RECT 2092.330 836.890 2093.510 838.070 ;
        RECT 2092.330 658.490 2093.510 659.670 ;
        RECT 2092.330 656.890 2093.510 658.070 ;
        RECT 2092.330 478.490 2093.510 479.670 ;
        RECT 2092.330 476.890 2093.510 478.070 ;
        RECT 2092.330 298.490 2093.510 299.670 ;
        RECT 2092.330 296.890 2093.510 298.070 ;
        RECT 2092.330 118.490 2093.510 119.670 ;
        RECT 2092.330 116.890 2093.510 118.070 ;
        RECT 2092.330 -16.710 2093.510 -15.530 ;
        RECT 2092.330 -18.310 2093.510 -17.130 ;
        RECT 2272.330 3536.810 2273.510 3537.990 ;
        RECT 2272.330 3535.210 2273.510 3536.390 ;
        RECT 2272.330 3358.490 2273.510 3359.670 ;
        RECT 2272.330 3356.890 2273.510 3358.070 ;
        RECT 2272.330 3178.490 2273.510 3179.670 ;
        RECT 2272.330 3176.890 2273.510 3178.070 ;
        RECT 2272.330 2998.490 2273.510 2999.670 ;
        RECT 2272.330 2996.890 2273.510 2998.070 ;
        RECT 2272.330 2818.490 2273.510 2819.670 ;
        RECT 2272.330 2816.890 2273.510 2818.070 ;
        RECT 2272.330 2638.490 2273.510 2639.670 ;
        RECT 2272.330 2636.890 2273.510 2638.070 ;
        RECT 2272.330 2458.490 2273.510 2459.670 ;
        RECT 2272.330 2456.890 2273.510 2458.070 ;
        RECT 2272.330 2278.490 2273.510 2279.670 ;
        RECT 2272.330 2276.890 2273.510 2278.070 ;
        RECT 2272.330 2098.490 2273.510 2099.670 ;
        RECT 2272.330 2096.890 2273.510 2098.070 ;
        RECT 2272.330 1918.490 2273.510 1919.670 ;
        RECT 2272.330 1916.890 2273.510 1918.070 ;
        RECT 2272.330 1738.490 2273.510 1739.670 ;
        RECT 2272.330 1736.890 2273.510 1738.070 ;
        RECT 2272.330 1558.490 2273.510 1559.670 ;
        RECT 2272.330 1556.890 2273.510 1558.070 ;
        RECT 2272.330 1378.490 2273.510 1379.670 ;
        RECT 2272.330 1376.890 2273.510 1378.070 ;
        RECT 2272.330 1198.490 2273.510 1199.670 ;
        RECT 2272.330 1196.890 2273.510 1198.070 ;
        RECT 2272.330 1018.490 2273.510 1019.670 ;
        RECT 2272.330 1016.890 2273.510 1018.070 ;
        RECT 2272.330 838.490 2273.510 839.670 ;
        RECT 2272.330 836.890 2273.510 838.070 ;
        RECT 2272.330 658.490 2273.510 659.670 ;
        RECT 2272.330 656.890 2273.510 658.070 ;
        RECT 2272.330 478.490 2273.510 479.670 ;
        RECT 2272.330 476.890 2273.510 478.070 ;
        RECT 2272.330 298.490 2273.510 299.670 ;
        RECT 2272.330 296.890 2273.510 298.070 ;
        RECT 2272.330 118.490 2273.510 119.670 ;
        RECT 2272.330 116.890 2273.510 118.070 ;
        RECT 2272.330 -16.710 2273.510 -15.530 ;
        RECT 2272.330 -18.310 2273.510 -17.130 ;
        RECT 2452.330 3536.810 2453.510 3537.990 ;
        RECT 2452.330 3535.210 2453.510 3536.390 ;
        RECT 2452.330 3358.490 2453.510 3359.670 ;
        RECT 2452.330 3356.890 2453.510 3358.070 ;
        RECT 2452.330 3178.490 2453.510 3179.670 ;
        RECT 2452.330 3176.890 2453.510 3178.070 ;
        RECT 2452.330 2998.490 2453.510 2999.670 ;
        RECT 2452.330 2996.890 2453.510 2998.070 ;
        RECT 2452.330 2818.490 2453.510 2819.670 ;
        RECT 2452.330 2816.890 2453.510 2818.070 ;
        RECT 2452.330 2638.490 2453.510 2639.670 ;
        RECT 2452.330 2636.890 2453.510 2638.070 ;
        RECT 2452.330 2458.490 2453.510 2459.670 ;
        RECT 2452.330 2456.890 2453.510 2458.070 ;
        RECT 2452.330 2278.490 2453.510 2279.670 ;
        RECT 2452.330 2276.890 2453.510 2278.070 ;
        RECT 2452.330 2098.490 2453.510 2099.670 ;
        RECT 2452.330 2096.890 2453.510 2098.070 ;
        RECT 2452.330 1918.490 2453.510 1919.670 ;
        RECT 2452.330 1916.890 2453.510 1918.070 ;
        RECT 2452.330 1738.490 2453.510 1739.670 ;
        RECT 2452.330 1736.890 2453.510 1738.070 ;
        RECT 2452.330 1558.490 2453.510 1559.670 ;
        RECT 2452.330 1556.890 2453.510 1558.070 ;
        RECT 2452.330 1378.490 2453.510 1379.670 ;
        RECT 2452.330 1376.890 2453.510 1378.070 ;
        RECT 2452.330 1198.490 2453.510 1199.670 ;
        RECT 2452.330 1196.890 2453.510 1198.070 ;
        RECT 2452.330 1018.490 2453.510 1019.670 ;
        RECT 2452.330 1016.890 2453.510 1018.070 ;
        RECT 2452.330 838.490 2453.510 839.670 ;
        RECT 2452.330 836.890 2453.510 838.070 ;
        RECT 2452.330 658.490 2453.510 659.670 ;
        RECT 2452.330 656.890 2453.510 658.070 ;
        RECT 2452.330 478.490 2453.510 479.670 ;
        RECT 2452.330 476.890 2453.510 478.070 ;
        RECT 2452.330 298.490 2453.510 299.670 ;
        RECT 2452.330 296.890 2453.510 298.070 ;
        RECT 2452.330 118.490 2453.510 119.670 ;
        RECT 2452.330 116.890 2453.510 118.070 ;
        RECT 2452.330 -16.710 2453.510 -15.530 ;
        RECT 2452.330 -18.310 2453.510 -17.130 ;
        RECT 2632.330 3536.810 2633.510 3537.990 ;
        RECT 2632.330 3535.210 2633.510 3536.390 ;
        RECT 2632.330 3358.490 2633.510 3359.670 ;
        RECT 2632.330 3356.890 2633.510 3358.070 ;
        RECT 2632.330 3178.490 2633.510 3179.670 ;
        RECT 2632.330 3176.890 2633.510 3178.070 ;
        RECT 2632.330 2998.490 2633.510 2999.670 ;
        RECT 2632.330 2996.890 2633.510 2998.070 ;
        RECT 2632.330 2818.490 2633.510 2819.670 ;
        RECT 2632.330 2816.890 2633.510 2818.070 ;
        RECT 2632.330 2638.490 2633.510 2639.670 ;
        RECT 2632.330 2636.890 2633.510 2638.070 ;
        RECT 2632.330 2458.490 2633.510 2459.670 ;
        RECT 2632.330 2456.890 2633.510 2458.070 ;
        RECT 2632.330 2278.490 2633.510 2279.670 ;
        RECT 2632.330 2276.890 2633.510 2278.070 ;
        RECT 2632.330 2098.490 2633.510 2099.670 ;
        RECT 2632.330 2096.890 2633.510 2098.070 ;
        RECT 2632.330 1918.490 2633.510 1919.670 ;
        RECT 2632.330 1916.890 2633.510 1918.070 ;
        RECT 2632.330 1738.490 2633.510 1739.670 ;
        RECT 2632.330 1736.890 2633.510 1738.070 ;
        RECT 2632.330 1558.490 2633.510 1559.670 ;
        RECT 2632.330 1556.890 2633.510 1558.070 ;
        RECT 2632.330 1378.490 2633.510 1379.670 ;
        RECT 2632.330 1376.890 2633.510 1378.070 ;
        RECT 2632.330 1198.490 2633.510 1199.670 ;
        RECT 2632.330 1196.890 2633.510 1198.070 ;
        RECT 2632.330 1018.490 2633.510 1019.670 ;
        RECT 2632.330 1016.890 2633.510 1018.070 ;
        RECT 2632.330 838.490 2633.510 839.670 ;
        RECT 2632.330 836.890 2633.510 838.070 ;
        RECT 2632.330 658.490 2633.510 659.670 ;
        RECT 2632.330 656.890 2633.510 658.070 ;
        RECT 2632.330 478.490 2633.510 479.670 ;
        RECT 2632.330 476.890 2633.510 478.070 ;
        RECT 2632.330 298.490 2633.510 299.670 ;
        RECT 2632.330 296.890 2633.510 298.070 ;
        RECT 2632.330 118.490 2633.510 119.670 ;
        RECT 2632.330 116.890 2633.510 118.070 ;
        RECT 2632.330 -16.710 2633.510 -15.530 ;
        RECT 2632.330 -18.310 2633.510 -17.130 ;
        RECT 2812.330 3536.810 2813.510 3537.990 ;
        RECT 2812.330 3535.210 2813.510 3536.390 ;
        RECT 2812.330 3358.490 2813.510 3359.670 ;
        RECT 2812.330 3356.890 2813.510 3358.070 ;
        RECT 2812.330 3178.490 2813.510 3179.670 ;
        RECT 2812.330 3176.890 2813.510 3178.070 ;
        RECT 2812.330 2998.490 2813.510 2999.670 ;
        RECT 2812.330 2996.890 2813.510 2998.070 ;
        RECT 2812.330 2818.490 2813.510 2819.670 ;
        RECT 2812.330 2816.890 2813.510 2818.070 ;
        RECT 2812.330 2638.490 2813.510 2639.670 ;
        RECT 2812.330 2636.890 2813.510 2638.070 ;
        RECT 2812.330 2458.490 2813.510 2459.670 ;
        RECT 2812.330 2456.890 2813.510 2458.070 ;
        RECT 2812.330 2278.490 2813.510 2279.670 ;
        RECT 2812.330 2276.890 2813.510 2278.070 ;
        RECT 2812.330 2098.490 2813.510 2099.670 ;
        RECT 2812.330 2096.890 2813.510 2098.070 ;
        RECT 2812.330 1918.490 2813.510 1919.670 ;
        RECT 2812.330 1916.890 2813.510 1918.070 ;
        RECT 2812.330 1738.490 2813.510 1739.670 ;
        RECT 2812.330 1736.890 2813.510 1738.070 ;
        RECT 2812.330 1558.490 2813.510 1559.670 ;
        RECT 2812.330 1556.890 2813.510 1558.070 ;
        RECT 2812.330 1378.490 2813.510 1379.670 ;
        RECT 2812.330 1376.890 2813.510 1378.070 ;
        RECT 2812.330 1198.490 2813.510 1199.670 ;
        RECT 2812.330 1196.890 2813.510 1198.070 ;
        RECT 2812.330 1018.490 2813.510 1019.670 ;
        RECT 2812.330 1016.890 2813.510 1018.070 ;
        RECT 2812.330 838.490 2813.510 839.670 ;
        RECT 2812.330 836.890 2813.510 838.070 ;
        RECT 2812.330 658.490 2813.510 659.670 ;
        RECT 2812.330 656.890 2813.510 658.070 ;
        RECT 2812.330 478.490 2813.510 479.670 ;
        RECT 2812.330 476.890 2813.510 478.070 ;
        RECT 2812.330 298.490 2813.510 299.670 ;
        RECT 2812.330 296.890 2813.510 298.070 ;
        RECT 2812.330 118.490 2813.510 119.670 ;
        RECT 2812.330 116.890 2813.510 118.070 ;
        RECT 2812.330 -16.710 2813.510 -15.530 ;
        RECT 2812.330 -18.310 2813.510 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3358.490 2942.490 3359.670 ;
        RECT 2941.310 3356.890 2942.490 3358.070 ;
        RECT 2941.310 3178.490 2942.490 3179.670 ;
        RECT 2941.310 3176.890 2942.490 3178.070 ;
        RECT 2941.310 2998.490 2942.490 2999.670 ;
        RECT 2941.310 2996.890 2942.490 2998.070 ;
        RECT 2941.310 2818.490 2942.490 2819.670 ;
        RECT 2941.310 2816.890 2942.490 2818.070 ;
        RECT 2941.310 2638.490 2942.490 2639.670 ;
        RECT 2941.310 2636.890 2942.490 2638.070 ;
        RECT 2941.310 2458.490 2942.490 2459.670 ;
        RECT 2941.310 2456.890 2942.490 2458.070 ;
        RECT 2941.310 2278.490 2942.490 2279.670 ;
        RECT 2941.310 2276.890 2942.490 2278.070 ;
        RECT 2941.310 2098.490 2942.490 2099.670 ;
        RECT 2941.310 2096.890 2942.490 2098.070 ;
        RECT 2941.310 1918.490 2942.490 1919.670 ;
        RECT 2941.310 1916.890 2942.490 1918.070 ;
        RECT 2941.310 1738.490 2942.490 1739.670 ;
        RECT 2941.310 1736.890 2942.490 1738.070 ;
        RECT 2941.310 1558.490 2942.490 1559.670 ;
        RECT 2941.310 1556.890 2942.490 1558.070 ;
        RECT 2941.310 1378.490 2942.490 1379.670 ;
        RECT 2941.310 1376.890 2942.490 1378.070 ;
        RECT 2941.310 1198.490 2942.490 1199.670 ;
        RECT 2941.310 1196.890 2942.490 1198.070 ;
        RECT 2941.310 1018.490 2942.490 1019.670 ;
        RECT 2941.310 1016.890 2942.490 1018.070 ;
        RECT 2941.310 838.490 2942.490 839.670 ;
        RECT 2941.310 836.890 2942.490 838.070 ;
        RECT 2941.310 658.490 2942.490 659.670 ;
        RECT 2941.310 656.890 2942.490 658.070 ;
        RECT 2941.310 478.490 2942.490 479.670 ;
        RECT 2941.310 476.890 2942.490 478.070 ;
        RECT 2941.310 298.490 2942.490 299.670 ;
        RECT 2941.310 296.890 2942.490 298.070 ;
        RECT 2941.310 118.490 2942.490 119.670 ;
        RECT 2941.310 116.890 2942.490 118.070 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.730 3538.050 -20.830 3538.110 ;
        RECT 111.470 3538.050 114.370 3538.110 ;
        RECT 291.470 3538.050 294.370 3538.110 ;
        RECT 471.470 3538.050 474.370 3538.110 ;
        RECT 651.470 3538.050 654.370 3538.110 ;
        RECT 831.470 3538.050 834.370 3538.110 ;
        RECT 1011.470 3538.050 1014.370 3538.110 ;
        RECT 1191.470 3538.050 1194.370 3538.110 ;
        RECT 1371.470 3538.050 1374.370 3538.110 ;
        RECT 1551.470 3538.050 1554.370 3538.110 ;
        RECT 1731.470 3538.050 1734.370 3538.110 ;
        RECT 1911.470 3538.050 1914.370 3538.110 ;
        RECT 2091.470 3538.050 2094.370 3538.110 ;
        RECT 2271.470 3538.050 2274.370 3538.110 ;
        RECT 2451.470 3538.050 2454.370 3538.110 ;
        RECT 2631.470 3538.050 2634.370 3538.110 ;
        RECT 2811.470 3538.050 2814.370 3538.110 ;
        RECT 2940.450 3538.050 2943.350 3538.110 ;
        RECT -23.730 3535.150 2943.350 3538.050 ;
        RECT -23.730 3535.090 -20.830 3535.150 ;
        RECT 111.470 3535.090 114.370 3535.150 ;
        RECT 291.470 3535.090 294.370 3535.150 ;
        RECT 471.470 3535.090 474.370 3535.150 ;
        RECT 651.470 3535.090 654.370 3535.150 ;
        RECT 831.470 3535.090 834.370 3535.150 ;
        RECT 1011.470 3535.090 1014.370 3535.150 ;
        RECT 1191.470 3535.090 1194.370 3535.150 ;
        RECT 1371.470 3535.090 1374.370 3535.150 ;
        RECT 1551.470 3535.090 1554.370 3535.150 ;
        RECT 1731.470 3535.090 1734.370 3535.150 ;
        RECT 1911.470 3535.090 1914.370 3535.150 ;
        RECT 2091.470 3535.090 2094.370 3535.150 ;
        RECT 2271.470 3535.090 2274.370 3535.150 ;
        RECT 2451.470 3535.090 2454.370 3535.150 ;
        RECT 2631.470 3535.090 2634.370 3535.150 ;
        RECT 2811.470 3535.090 2814.370 3535.150 ;
        RECT 2940.450 3535.090 2943.350 3535.150 ;
        RECT -23.730 3359.730 -20.830 3359.790 ;
        RECT 111.470 3359.730 114.370 3359.790 ;
        RECT 291.470 3359.730 294.370 3359.790 ;
        RECT 471.470 3359.730 474.370 3359.790 ;
        RECT 651.470 3359.730 654.370 3359.790 ;
        RECT 831.470 3359.730 834.370 3359.790 ;
        RECT 1011.470 3359.730 1014.370 3359.790 ;
        RECT 1191.470 3359.730 1194.370 3359.790 ;
        RECT 1371.470 3359.730 1374.370 3359.790 ;
        RECT 1551.470 3359.730 1554.370 3359.790 ;
        RECT 1731.470 3359.730 1734.370 3359.790 ;
        RECT 1911.470 3359.730 1914.370 3359.790 ;
        RECT 2091.470 3359.730 2094.370 3359.790 ;
        RECT 2271.470 3359.730 2274.370 3359.790 ;
        RECT 2451.470 3359.730 2454.370 3359.790 ;
        RECT 2631.470 3359.730 2634.370 3359.790 ;
        RECT 2811.470 3359.730 2814.370 3359.790 ;
        RECT 2940.450 3359.730 2943.350 3359.790 ;
        RECT -23.730 3356.830 2943.350 3359.730 ;
        RECT -23.730 3356.770 -20.830 3356.830 ;
        RECT 111.470 3356.770 114.370 3356.830 ;
        RECT 291.470 3356.770 294.370 3356.830 ;
        RECT 471.470 3356.770 474.370 3356.830 ;
        RECT 651.470 3356.770 654.370 3356.830 ;
        RECT 831.470 3356.770 834.370 3356.830 ;
        RECT 1011.470 3356.770 1014.370 3356.830 ;
        RECT 1191.470 3356.770 1194.370 3356.830 ;
        RECT 1371.470 3356.770 1374.370 3356.830 ;
        RECT 1551.470 3356.770 1554.370 3356.830 ;
        RECT 1731.470 3356.770 1734.370 3356.830 ;
        RECT 1911.470 3356.770 1914.370 3356.830 ;
        RECT 2091.470 3356.770 2094.370 3356.830 ;
        RECT 2271.470 3356.770 2274.370 3356.830 ;
        RECT 2451.470 3356.770 2454.370 3356.830 ;
        RECT 2631.470 3356.770 2634.370 3356.830 ;
        RECT 2811.470 3356.770 2814.370 3356.830 ;
        RECT 2940.450 3356.770 2943.350 3356.830 ;
        RECT -23.730 3179.730 -20.830 3179.790 ;
        RECT 111.470 3179.730 114.370 3179.790 ;
        RECT 291.470 3179.730 294.370 3179.790 ;
        RECT 471.470 3179.730 474.370 3179.790 ;
        RECT 651.470 3179.730 654.370 3179.790 ;
        RECT 831.470 3179.730 834.370 3179.790 ;
        RECT 1011.470 3179.730 1014.370 3179.790 ;
        RECT 1191.470 3179.730 1194.370 3179.790 ;
        RECT 1371.470 3179.730 1374.370 3179.790 ;
        RECT 1551.470 3179.730 1554.370 3179.790 ;
        RECT 1731.470 3179.730 1734.370 3179.790 ;
        RECT 1911.470 3179.730 1914.370 3179.790 ;
        RECT 2091.470 3179.730 2094.370 3179.790 ;
        RECT 2271.470 3179.730 2274.370 3179.790 ;
        RECT 2451.470 3179.730 2454.370 3179.790 ;
        RECT 2631.470 3179.730 2634.370 3179.790 ;
        RECT 2811.470 3179.730 2814.370 3179.790 ;
        RECT 2940.450 3179.730 2943.350 3179.790 ;
        RECT -23.730 3176.830 2943.350 3179.730 ;
        RECT -23.730 3176.770 -20.830 3176.830 ;
        RECT 111.470 3176.770 114.370 3176.830 ;
        RECT 291.470 3176.770 294.370 3176.830 ;
        RECT 471.470 3176.770 474.370 3176.830 ;
        RECT 651.470 3176.770 654.370 3176.830 ;
        RECT 831.470 3176.770 834.370 3176.830 ;
        RECT 1011.470 3176.770 1014.370 3176.830 ;
        RECT 1191.470 3176.770 1194.370 3176.830 ;
        RECT 1371.470 3176.770 1374.370 3176.830 ;
        RECT 1551.470 3176.770 1554.370 3176.830 ;
        RECT 1731.470 3176.770 1734.370 3176.830 ;
        RECT 1911.470 3176.770 1914.370 3176.830 ;
        RECT 2091.470 3176.770 2094.370 3176.830 ;
        RECT 2271.470 3176.770 2274.370 3176.830 ;
        RECT 2451.470 3176.770 2454.370 3176.830 ;
        RECT 2631.470 3176.770 2634.370 3176.830 ;
        RECT 2811.470 3176.770 2814.370 3176.830 ;
        RECT 2940.450 3176.770 2943.350 3176.830 ;
        RECT -23.730 2999.730 -20.830 2999.790 ;
        RECT 111.470 2999.730 114.370 2999.790 ;
        RECT 291.470 2999.730 294.370 2999.790 ;
        RECT 471.470 2999.730 474.370 2999.790 ;
        RECT 651.470 2999.730 654.370 2999.790 ;
        RECT 831.470 2999.730 834.370 2999.790 ;
        RECT 1011.470 2999.730 1014.370 2999.790 ;
        RECT 1191.470 2999.730 1194.370 2999.790 ;
        RECT 1371.470 2999.730 1374.370 2999.790 ;
        RECT 1551.470 2999.730 1554.370 2999.790 ;
        RECT 1731.470 2999.730 1734.370 2999.790 ;
        RECT 1911.470 2999.730 1914.370 2999.790 ;
        RECT 2091.470 2999.730 2094.370 2999.790 ;
        RECT 2271.470 2999.730 2274.370 2999.790 ;
        RECT 2451.470 2999.730 2454.370 2999.790 ;
        RECT 2631.470 2999.730 2634.370 2999.790 ;
        RECT 2811.470 2999.730 2814.370 2999.790 ;
        RECT 2940.450 2999.730 2943.350 2999.790 ;
        RECT -23.730 2996.830 2943.350 2999.730 ;
        RECT -23.730 2996.770 -20.830 2996.830 ;
        RECT 111.470 2996.770 114.370 2996.830 ;
        RECT 291.470 2996.770 294.370 2996.830 ;
        RECT 471.470 2996.770 474.370 2996.830 ;
        RECT 651.470 2996.770 654.370 2996.830 ;
        RECT 831.470 2996.770 834.370 2996.830 ;
        RECT 1011.470 2996.770 1014.370 2996.830 ;
        RECT 1191.470 2996.770 1194.370 2996.830 ;
        RECT 1371.470 2996.770 1374.370 2996.830 ;
        RECT 1551.470 2996.770 1554.370 2996.830 ;
        RECT 1731.470 2996.770 1734.370 2996.830 ;
        RECT 1911.470 2996.770 1914.370 2996.830 ;
        RECT 2091.470 2996.770 2094.370 2996.830 ;
        RECT 2271.470 2996.770 2274.370 2996.830 ;
        RECT 2451.470 2996.770 2454.370 2996.830 ;
        RECT 2631.470 2996.770 2634.370 2996.830 ;
        RECT 2811.470 2996.770 2814.370 2996.830 ;
        RECT 2940.450 2996.770 2943.350 2996.830 ;
        RECT -23.730 2819.730 -20.830 2819.790 ;
        RECT 111.470 2819.730 114.370 2819.790 ;
        RECT 291.470 2819.730 294.370 2819.790 ;
        RECT 471.470 2819.730 474.370 2819.790 ;
        RECT 651.470 2819.730 654.370 2819.790 ;
        RECT 831.470 2819.730 834.370 2819.790 ;
        RECT 1011.470 2819.730 1014.370 2819.790 ;
        RECT 1191.470 2819.730 1194.370 2819.790 ;
        RECT 1371.470 2819.730 1374.370 2819.790 ;
        RECT 1551.470 2819.730 1554.370 2819.790 ;
        RECT 1731.470 2819.730 1734.370 2819.790 ;
        RECT 1911.470 2819.730 1914.370 2819.790 ;
        RECT 2091.470 2819.730 2094.370 2819.790 ;
        RECT 2271.470 2819.730 2274.370 2819.790 ;
        RECT 2451.470 2819.730 2454.370 2819.790 ;
        RECT 2631.470 2819.730 2634.370 2819.790 ;
        RECT 2811.470 2819.730 2814.370 2819.790 ;
        RECT 2940.450 2819.730 2943.350 2819.790 ;
        RECT -23.730 2816.830 2943.350 2819.730 ;
        RECT -23.730 2816.770 -20.830 2816.830 ;
        RECT 111.470 2816.770 114.370 2816.830 ;
        RECT 291.470 2816.770 294.370 2816.830 ;
        RECT 471.470 2816.770 474.370 2816.830 ;
        RECT 651.470 2816.770 654.370 2816.830 ;
        RECT 831.470 2816.770 834.370 2816.830 ;
        RECT 1011.470 2816.770 1014.370 2816.830 ;
        RECT 1191.470 2816.770 1194.370 2816.830 ;
        RECT 1371.470 2816.770 1374.370 2816.830 ;
        RECT 1551.470 2816.770 1554.370 2816.830 ;
        RECT 1731.470 2816.770 1734.370 2816.830 ;
        RECT 1911.470 2816.770 1914.370 2816.830 ;
        RECT 2091.470 2816.770 2094.370 2816.830 ;
        RECT 2271.470 2816.770 2274.370 2816.830 ;
        RECT 2451.470 2816.770 2454.370 2816.830 ;
        RECT 2631.470 2816.770 2634.370 2816.830 ;
        RECT 2811.470 2816.770 2814.370 2816.830 ;
        RECT 2940.450 2816.770 2943.350 2816.830 ;
        RECT -23.730 2639.730 -20.830 2639.790 ;
        RECT 111.470 2639.730 114.370 2639.790 ;
        RECT 291.470 2639.730 294.370 2639.790 ;
        RECT 471.470 2639.730 474.370 2639.790 ;
        RECT 651.470 2639.730 654.370 2639.790 ;
        RECT 831.470 2639.730 834.370 2639.790 ;
        RECT 1011.470 2639.730 1014.370 2639.790 ;
        RECT 1191.470 2639.730 1194.370 2639.790 ;
        RECT 1371.470 2639.730 1374.370 2639.790 ;
        RECT 1551.470 2639.730 1554.370 2639.790 ;
        RECT 1731.470 2639.730 1734.370 2639.790 ;
        RECT 1911.470 2639.730 1914.370 2639.790 ;
        RECT 2091.470 2639.730 2094.370 2639.790 ;
        RECT 2271.470 2639.730 2274.370 2639.790 ;
        RECT 2451.470 2639.730 2454.370 2639.790 ;
        RECT 2631.470 2639.730 2634.370 2639.790 ;
        RECT 2811.470 2639.730 2814.370 2639.790 ;
        RECT 2940.450 2639.730 2943.350 2639.790 ;
        RECT -23.730 2636.830 2943.350 2639.730 ;
        RECT -23.730 2636.770 -20.830 2636.830 ;
        RECT 111.470 2636.770 114.370 2636.830 ;
        RECT 291.470 2636.770 294.370 2636.830 ;
        RECT 471.470 2636.770 474.370 2636.830 ;
        RECT 651.470 2636.770 654.370 2636.830 ;
        RECT 831.470 2636.770 834.370 2636.830 ;
        RECT 1011.470 2636.770 1014.370 2636.830 ;
        RECT 1191.470 2636.770 1194.370 2636.830 ;
        RECT 1371.470 2636.770 1374.370 2636.830 ;
        RECT 1551.470 2636.770 1554.370 2636.830 ;
        RECT 1731.470 2636.770 1734.370 2636.830 ;
        RECT 1911.470 2636.770 1914.370 2636.830 ;
        RECT 2091.470 2636.770 2094.370 2636.830 ;
        RECT 2271.470 2636.770 2274.370 2636.830 ;
        RECT 2451.470 2636.770 2454.370 2636.830 ;
        RECT 2631.470 2636.770 2634.370 2636.830 ;
        RECT 2811.470 2636.770 2814.370 2636.830 ;
        RECT 2940.450 2636.770 2943.350 2636.830 ;
        RECT -23.730 2459.730 -20.830 2459.790 ;
        RECT 111.470 2459.730 114.370 2459.790 ;
        RECT 291.470 2459.730 294.370 2459.790 ;
        RECT 471.470 2459.730 474.370 2459.790 ;
        RECT 651.470 2459.730 654.370 2459.790 ;
        RECT 831.470 2459.730 834.370 2459.790 ;
        RECT 1011.470 2459.730 1014.370 2459.790 ;
        RECT 1191.470 2459.730 1194.370 2459.790 ;
        RECT 1371.470 2459.730 1374.370 2459.790 ;
        RECT 1551.470 2459.730 1554.370 2459.790 ;
        RECT 1731.470 2459.730 1734.370 2459.790 ;
        RECT 1911.470 2459.730 1914.370 2459.790 ;
        RECT 2091.470 2459.730 2094.370 2459.790 ;
        RECT 2271.470 2459.730 2274.370 2459.790 ;
        RECT 2451.470 2459.730 2454.370 2459.790 ;
        RECT 2631.470 2459.730 2634.370 2459.790 ;
        RECT 2811.470 2459.730 2814.370 2459.790 ;
        RECT 2940.450 2459.730 2943.350 2459.790 ;
        RECT -23.730 2456.830 2943.350 2459.730 ;
        RECT -23.730 2456.770 -20.830 2456.830 ;
        RECT 111.470 2456.770 114.370 2456.830 ;
        RECT 291.470 2456.770 294.370 2456.830 ;
        RECT 471.470 2456.770 474.370 2456.830 ;
        RECT 651.470 2456.770 654.370 2456.830 ;
        RECT 831.470 2456.770 834.370 2456.830 ;
        RECT 1011.470 2456.770 1014.370 2456.830 ;
        RECT 1191.470 2456.770 1194.370 2456.830 ;
        RECT 1371.470 2456.770 1374.370 2456.830 ;
        RECT 1551.470 2456.770 1554.370 2456.830 ;
        RECT 1731.470 2456.770 1734.370 2456.830 ;
        RECT 1911.470 2456.770 1914.370 2456.830 ;
        RECT 2091.470 2456.770 2094.370 2456.830 ;
        RECT 2271.470 2456.770 2274.370 2456.830 ;
        RECT 2451.470 2456.770 2454.370 2456.830 ;
        RECT 2631.470 2456.770 2634.370 2456.830 ;
        RECT 2811.470 2456.770 2814.370 2456.830 ;
        RECT 2940.450 2456.770 2943.350 2456.830 ;
        RECT -23.730 2279.730 -20.830 2279.790 ;
        RECT 111.470 2279.730 114.370 2279.790 ;
        RECT 291.470 2279.730 294.370 2279.790 ;
        RECT 471.470 2279.730 474.370 2279.790 ;
        RECT 651.470 2279.730 654.370 2279.790 ;
        RECT 831.470 2279.730 834.370 2279.790 ;
        RECT 1011.470 2279.730 1014.370 2279.790 ;
        RECT 1191.470 2279.730 1194.370 2279.790 ;
        RECT 1371.470 2279.730 1374.370 2279.790 ;
        RECT 1551.470 2279.730 1554.370 2279.790 ;
        RECT 1731.470 2279.730 1734.370 2279.790 ;
        RECT 1911.470 2279.730 1914.370 2279.790 ;
        RECT 2091.470 2279.730 2094.370 2279.790 ;
        RECT 2271.470 2279.730 2274.370 2279.790 ;
        RECT 2451.470 2279.730 2454.370 2279.790 ;
        RECT 2631.470 2279.730 2634.370 2279.790 ;
        RECT 2811.470 2279.730 2814.370 2279.790 ;
        RECT 2940.450 2279.730 2943.350 2279.790 ;
        RECT -23.730 2276.830 2943.350 2279.730 ;
        RECT -23.730 2276.770 -20.830 2276.830 ;
        RECT 111.470 2276.770 114.370 2276.830 ;
        RECT 291.470 2276.770 294.370 2276.830 ;
        RECT 471.470 2276.770 474.370 2276.830 ;
        RECT 651.470 2276.770 654.370 2276.830 ;
        RECT 831.470 2276.770 834.370 2276.830 ;
        RECT 1011.470 2276.770 1014.370 2276.830 ;
        RECT 1191.470 2276.770 1194.370 2276.830 ;
        RECT 1371.470 2276.770 1374.370 2276.830 ;
        RECT 1551.470 2276.770 1554.370 2276.830 ;
        RECT 1731.470 2276.770 1734.370 2276.830 ;
        RECT 1911.470 2276.770 1914.370 2276.830 ;
        RECT 2091.470 2276.770 2094.370 2276.830 ;
        RECT 2271.470 2276.770 2274.370 2276.830 ;
        RECT 2451.470 2276.770 2454.370 2276.830 ;
        RECT 2631.470 2276.770 2634.370 2276.830 ;
        RECT 2811.470 2276.770 2814.370 2276.830 ;
        RECT 2940.450 2276.770 2943.350 2276.830 ;
        RECT -23.730 2099.730 -20.830 2099.790 ;
        RECT 111.470 2099.730 114.370 2099.790 ;
        RECT 291.470 2099.730 294.370 2099.790 ;
        RECT 471.470 2099.730 474.370 2099.790 ;
        RECT 651.470 2099.730 654.370 2099.790 ;
        RECT 831.470 2099.730 834.370 2099.790 ;
        RECT 1011.470 2099.730 1014.370 2099.790 ;
        RECT 1191.470 2099.730 1194.370 2099.790 ;
        RECT 1371.470 2099.730 1374.370 2099.790 ;
        RECT 1551.470 2099.730 1554.370 2099.790 ;
        RECT 1731.470 2099.730 1734.370 2099.790 ;
        RECT 1911.470 2099.730 1914.370 2099.790 ;
        RECT 2091.470 2099.730 2094.370 2099.790 ;
        RECT 2271.470 2099.730 2274.370 2099.790 ;
        RECT 2451.470 2099.730 2454.370 2099.790 ;
        RECT 2631.470 2099.730 2634.370 2099.790 ;
        RECT 2811.470 2099.730 2814.370 2099.790 ;
        RECT 2940.450 2099.730 2943.350 2099.790 ;
        RECT -23.730 2096.830 2943.350 2099.730 ;
        RECT -23.730 2096.770 -20.830 2096.830 ;
        RECT 111.470 2096.770 114.370 2096.830 ;
        RECT 291.470 2096.770 294.370 2096.830 ;
        RECT 471.470 2096.770 474.370 2096.830 ;
        RECT 651.470 2096.770 654.370 2096.830 ;
        RECT 831.470 2096.770 834.370 2096.830 ;
        RECT 1011.470 2096.770 1014.370 2096.830 ;
        RECT 1191.470 2096.770 1194.370 2096.830 ;
        RECT 1371.470 2096.770 1374.370 2096.830 ;
        RECT 1551.470 2096.770 1554.370 2096.830 ;
        RECT 1731.470 2096.770 1734.370 2096.830 ;
        RECT 1911.470 2096.770 1914.370 2096.830 ;
        RECT 2091.470 2096.770 2094.370 2096.830 ;
        RECT 2271.470 2096.770 2274.370 2096.830 ;
        RECT 2451.470 2096.770 2454.370 2096.830 ;
        RECT 2631.470 2096.770 2634.370 2096.830 ;
        RECT 2811.470 2096.770 2814.370 2096.830 ;
        RECT 2940.450 2096.770 2943.350 2096.830 ;
        RECT -23.730 1919.730 -20.830 1919.790 ;
        RECT 111.470 1919.730 114.370 1919.790 ;
        RECT 291.470 1919.730 294.370 1919.790 ;
        RECT 471.470 1919.730 474.370 1919.790 ;
        RECT 651.470 1919.730 654.370 1919.790 ;
        RECT 831.470 1919.730 834.370 1919.790 ;
        RECT 1011.470 1919.730 1014.370 1919.790 ;
        RECT 1191.470 1919.730 1194.370 1919.790 ;
        RECT 1371.470 1919.730 1374.370 1919.790 ;
        RECT 1551.470 1919.730 1554.370 1919.790 ;
        RECT 1731.470 1919.730 1734.370 1919.790 ;
        RECT 1911.470 1919.730 1914.370 1919.790 ;
        RECT 2091.470 1919.730 2094.370 1919.790 ;
        RECT 2271.470 1919.730 2274.370 1919.790 ;
        RECT 2451.470 1919.730 2454.370 1919.790 ;
        RECT 2631.470 1919.730 2634.370 1919.790 ;
        RECT 2811.470 1919.730 2814.370 1919.790 ;
        RECT 2940.450 1919.730 2943.350 1919.790 ;
        RECT -23.730 1916.830 2943.350 1919.730 ;
        RECT -23.730 1916.770 -20.830 1916.830 ;
        RECT 111.470 1916.770 114.370 1916.830 ;
        RECT 291.470 1916.770 294.370 1916.830 ;
        RECT 471.470 1916.770 474.370 1916.830 ;
        RECT 651.470 1916.770 654.370 1916.830 ;
        RECT 831.470 1916.770 834.370 1916.830 ;
        RECT 1011.470 1916.770 1014.370 1916.830 ;
        RECT 1191.470 1916.770 1194.370 1916.830 ;
        RECT 1371.470 1916.770 1374.370 1916.830 ;
        RECT 1551.470 1916.770 1554.370 1916.830 ;
        RECT 1731.470 1916.770 1734.370 1916.830 ;
        RECT 1911.470 1916.770 1914.370 1916.830 ;
        RECT 2091.470 1916.770 2094.370 1916.830 ;
        RECT 2271.470 1916.770 2274.370 1916.830 ;
        RECT 2451.470 1916.770 2454.370 1916.830 ;
        RECT 2631.470 1916.770 2634.370 1916.830 ;
        RECT 2811.470 1916.770 2814.370 1916.830 ;
        RECT 2940.450 1916.770 2943.350 1916.830 ;
        RECT -23.730 1739.730 -20.830 1739.790 ;
        RECT 111.470 1739.730 114.370 1739.790 ;
        RECT 291.470 1739.730 294.370 1739.790 ;
        RECT 471.470 1739.730 474.370 1739.790 ;
        RECT 651.470 1739.730 654.370 1739.790 ;
        RECT 831.470 1739.730 834.370 1739.790 ;
        RECT 1011.470 1739.730 1014.370 1739.790 ;
        RECT 1191.470 1739.730 1194.370 1739.790 ;
        RECT 1371.470 1739.730 1374.370 1739.790 ;
        RECT 1551.470 1739.730 1554.370 1739.790 ;
        RECT 1731.470 1739.730 1734.370 1739.790 ;
        RECT 1911.470 1739.730 1914.370 1739.790 ;
        RECT 2091.470 1739.730 2094.370 1739.790 ;
        RECT 2271.470 1739.730 2274.370 1739.790 ;
        RECT 2451.470 1739.730 2454.370 1739.790 ;
        RECT 2631.470 1739.730 2634.370 1739.790 ;
        RECT 2811.470 1739.730 2814.370 1739.790 ;
        RECT 2940.450 1739.730 2943.350 1739.790 ;
        RECT -23.730 1736.830 2943.350 1739.730 ;
        RECT -23.730 1736.770 -20.830 1736.830 ;
        RECT 111.470 1736.770 114.370 1736.830 ;
        RECT 291.470 1736.770 294.370 1736.830 ;
        RECT 471.470 1736.770 474.370 1736.830 ;
        RECT 651.470 1736.770 654.370 1736.830 ;
        RECT 831.470 1736.770 834.370 1736.830 ;
        RECT 1011.470 1736.770 1014.370 1736.830 ;
        RECT 1191.470 1736.770 1194.370 1736.830 ;
        RECT 1371.470 1736.770 1374.370 1736.830 ;
        RECT 1551.470 1736.770 1554.370 1736.830 ;
        RECT 1731.470 1736.770 1734.370 1736.830 ;
        RECT 1911.470 1736.770 1914.370 1736.830 ;
        RECT 2091.470 1736.770 2094.370 1736.830 ;
        RECT 2271.470 1736.770 2274.370 1736.830 ;
        RECT 2451.470 1736.770 2454.370 1736.830 ;
        RECT 2631.470 1736.770 2634.370 1736.830 ;
        RECT 2811.470 1736.770 2814.370 1736.830 ;
        RECT 2940.450 1736.770 2943.350 1736.830 ;
        RECT -23.730 1559.730 -20.830 1559.790 ;
        RECT 111.470 1559.730 114.370 1559.790 ;
        RECT 291.470 1559.730 294.370 1559.790 ;
        RECT 471.470 1559.730 474.370 1559.790 ;
        RECT 651.470 1559.730 654.370 1559.790 ;
        RECT 831.470 1559.730 834.370 1559.790 ;
        RECT 1011.470 1559.730 1014.370 1559.790 ;
        RECT 1191.470 1559.730 1194.370 1559.790 ;
        RECT 1371.470 1559.730 1374.370 1559.790 ;
        RECT 1551.470 1559.730 1554.370 1559.790 ;
        RECT 1731.470 1559.730 1734.370 1559.790 ;
        RECT 1911.470 1559.730 1914.370 1559.790 ;
        RECT 2091.470 1559.730 2094.370 1559.790 ;
        RECT 2271.470 1559.730 2274.370 1559.790 ;
        RECT 2451.470 1559.730 2454.370 1559.790 ;
        RECT 2631.470 1559.730 2634.370 1559.790 ;
        RECT 2811.470 1559.730 2814.370 1559.790 ;
        RECT 2940.450 1559.730 2943.350 1559.790 ;
        RECT -23.730 1556.830 2943.350 1559.730 ;
        RECT -23.730 1556.770 -20.830 1556.830 ;
        RECT 111.470 1556.770 114.370 1556.830 ;
        RECT 291.470 1556.770 294.370 1556.830 ;
        RECT 471.470 1556.770 474.370 1556.830 ;
        RECT 651.470 1556.770 654.370 1556.830 ;
        RECT 831.470 1556.770 834.370 1556.830 ;
        RECT 1011.470 1556.770 1014.370 1556.830 ;
        RECT 1191.470 1556.770 1194.370 1556.830 ;
        RECT 1371.470 1556.770 1374.370 1556.830 ;
        RECT 1551.470 1556.770 1554.370 1556.830 ;
        RECT 1731.470 1556.770 1734.370 1556.830 ;
        RECT 1911.470 1556.770 1914.370 1556.830 ;
        RECT 2091.470 1556.770 2094.370 1556.830 ;
        RECT 2271.470 1556.770 2274.370 1556.830 ;
        RECT 2451.470 1556.770 2454.370 1556.830 ;
        RECT 2631.470 1556.770 2634.370 1556.830 ;
        RECT 2811.470 1556.770 2814.370 1556.830 ;
        RECT 2940.450 1556.770 2943.350 1556.830 ;
        RECT -23.730 1379.730 -20.830 1379.790 ;
        RECT 111.470 1379.730 114.370 1379.790 ;
        RECT 291.470 1379.730 294.370 1379.790 ;
        RECT 471.470 1379.730 474.370 1379.790 ;
        RECT 651.470 1379.730 654.370 1379.790 ;
        RECT 831.470 1379.730 834.370 1379.790 ;
        RECT 1011.470 1379.730 1014.370 1379.790 ;
        RECT 1191.470 1379.730 1194.370 1379.790 ;
        RECT 1371.470 1379.730 1374.370 1379.790 ;
        RECT 1551.470 1379.730 1554.370 1379.790 ;
        RECT 1731.470 1379.730 1734.370 1379.790 ;
        RECT 1911.470 1379.730 1914.370 1379.790 ;
        RECT 2091.470 1379.730 2094.370 1379.790 ;
        RECT 2271.470 1379.730 2274.370 1379.790 ;
        RECT 2451.470 1379.730 2454.370 1379.790 ;
        RECT 2631.470 1379.730 2634.370 1379.790 ;
        RECT 2811.470 1379.730 2814.370 1379.790 ;
        RECT 2940.450 1379.730 2943.350 1379.790 ;
        RECT -23.730 1376.830 2943.350 1379.730 ;
        RECT -23.730 1376.770 -20.830 1376.830 ;
        RECT 111.470 1376.770 114.370 1376.830 ;
        RECT 291.470 1376.770 294.370 1376.830 ;
        RECT 471.470 1376.770 474.370 1376.830 ;
        RECT 651.470 1376.770 654.370 1376.830 ;
        RECT 831.470 1376.770 834.370 1376.830 ;
        RECT 1011.470 1376.770 1014.370 1376.830 ;
        RECT 1191.470 1376.770 1194.370 1376.830 ;
        RECT 1371.470 1376.770 1374.370 1376.830 ;
        RECT 1551.470 1376.770 1554.370 1376.830 ;
        RECT 1731.470 1376.770 1734.370 1376.830 ;
        RECT 1911.470 1376.770 1914.370 1376.830 ;
        RECT 2091.470 1376.770 2094.370 1376.830 ;
        RECT 2271.470 1376.770 2274.370 1376.830 ;
        RECT 2451.470 1376.770 2454.370 1376.830 ;
        RECT 2631.470 1376.770 2634.370 1376.830 ;
        RECT 2811.470 1376.770 2814.370 1376.830 ;
        RECT 2940.450 1376.770 2943.350 1376.830 ;
        RECT -23.730 1199.730 -20.830 1199.790 ;
        RECT 111.470 1199.730 114.370 1199.790 ;
        RECT 291.470 1199.730 294.370 1199.790 ;
        RECT 471.470 1199.730 474.370 1199.790 ;
        RECT 651.470 1199.730 654.370 1199.790 ;
        RECT 831.470 1199.730 834.370 1199.790 ;
        RECT 1011.470 1199.730 1014.370 1199.790 ;
        RECT 1191.470 1199.730 1194.370 1199.790 ;
        RECT 1371.470 1199.730 1374.370 1199.790 ;
        RECT 1551.470 1199.730 1554.370 1199.790 ;
        RECT 1731.470 1199.730 1734.370 1199.790 ;
        RECT 1911.470 1199.730 1914.370 1199.790 ;
        RECT 2091.470 1199.730 2094.370 1199.790 ;
        RECT 2271.470 1199.730 2274.370 1199.790 ;
        RECT 2451.470 1199.730 2454.370 1199.790 ;
        RECT 2631.470 1199.730 2634.370 1199.790 ;
        RECT 2811.470 1199.730 2814.370 1199.790 ;
        RECT 2940.450 1199.730 2943.350 1199.790 ;
        RECT -23.730 1196.830 2943.350 1199.730 ;
        RECT -23.730 1196.770 -20.830 1196.830 ;
        RECT 111.470 1196.770 114.370 1196.830 ;
        RECT 291.470 1196.770 294.370 1196.830 ;
        RECT 471.470 1196.770 474.370 1196.830 ;
        RECT 651.470 1196.770 654.370 1196.830 ;
        RECT 831.470 1196.770 834.370 1196.830 ;
        RECT 1011.470 1196.770 1014.370 1196.830 ;
        RECT 1191.470 1196.770 1194.370 1196.830 ;
        RECT 1371.470 1196.770 1374.370 1196.830 ;
        RECT 1551.470 1196.770 1554.370 1196.830 ;
        RECT 1731.470 1196.770 1734.370 1196.830 ;
        RECT 1911.470 1196.770 1914.370 1196.830 ;
        RECT 2091.470 1196.770 2094.370 1196.830 ;
        RECT 2271.470 1196.770 2274.370 1196.830 ;
        RECT 2451.470 1196.770 2454.370 1196.830 ;
        RECT 2631.470 1196.770 2634.370 1196.830 ;
        RECT 2811.470 1196.770 2814.370 1196.830 ;
        RECT 2940.450 1196.770 2943.350 1196.830 ;
        RECT -23.730 1019.730 -20.830 1019.790 ;
        RECT 111.470 1019.730 114.370 1019.790 ;
        RECT 291.470 1019.730 294.370 1019.790 ;
        RECT 471.470 1019.730 474.370 1019.790 ;
        RECT 651.470 1019.730 654.370 1019.790 ;
        RECT 831.470 1019.730 834.370 1019.790 ;
        RECT 1011.470 1019.730 1014.370 1019.790 ;
        RECT 1191.470 1019.730 1194.370 1019.790 ;
        RECT 1371.470 1019.730 1374.370 1019.790 ;
        RECT 1551.470 1019.730 1554.370 1019.790 ;
        RECT 1731.470 1019.730 1734.370 1019.790 ;
        RECT 1911.470 1019.730 1914.370 1019.790 ;
        RECT 2091.470 1019.730 2094.370 1019.790 ;
        RECT 2271.470 1019.730 2274.370 1019.790 ;
        RECT 2451.470 1019.730 2454.370 1019.790 ;
        RECT 2631.470 1019.730 2634.370 1019.790 ;
        RECT 2811.470 1019.730 2814.370 1019.790 ;
        RECT 2940.450 1019.730 2943.350 1019.790 ;
        RECT -23.730 1016.830 2943.350 1019.730 ;
        RECT -23.730 1016.770 -20.830 1016.830 ;
        RECT 111.470 1016.770 114.370 1016.830 ;
        RECT 291.470 1016.770 294.370 1016.830 ;
        RECT 471.470 1016.770 474.370 1016.830 ;
        RECT 651.470 1016.770 654.370 1016.830 ;
        RECT 831.470 1016.770 834.370 1016.830 ;
        RECT 1011.470 1016.770 1014.370 1016.830 ;
        RECT 1191.470 1016.770 1194.370 1016.830 ;
        RECT 1371.470 1016.770 1374.370 1016.830 ;
        RECT 1551.470 1016.770 1554.370 1016.830 ;
        RECT 1731.470 1016.770 1734.370 1016.830 ;
        RECT 1911.470 1016.770 1914.370 1016.830 ;
        RECT 2091.470 1016.770 2094.370 1016.830 ;
        RECT 2271.470 1016.770 2274.370 1016.830 ;
        RECT 2451.470 1016.770 2454.370 1016.830 ;
        RECT 2631.470 1016.770 2634.370 1016.830 ;
        RECT 2811.470 1016.770 2814.370 1016.830 ;
        RECT 2940.450 1016.770 2943.350 1016.830 ;
        RECT -23.730 839.730 -20.830 839.790 ;
        RECT 111.470 839.730 114.370 839.790 ;
        RECT 291.470 839.730 294.370 839.790 ;
        RECT 471.470 839.730 474.370 839.790 ;
        RECT 651.470 839.730 654.370 839.790 ;
        RECT 831.470 839.730 834.370 839.790 ;
        RECT 1011.470 839.730 1014.370 839.790 ;
        RECT 1191.470 839.730 1194.370 839.790 ;
        RECT 1371.470 839.730 1374.370 839.790 ;
        RECT 1551.470 839.730 1554.370 839.790 ;
        RECT 1731.470 839.730 1734.370 839.790 ;
        RECT 1911.470 839.730 1914.370 839.790 ;
        RECT 2091.470 839.730 2094.370 839.790 ;
        RECT 2271.470 839.730 2274.370 839.790 ;
        RECT 2451.470 839.730 2454.370 839.790 ;
        RECT 2631.470 839.730 2634.370 839.790 ;
        RECT 2811.470 839.730 2814.370 839.790 ;
        RECT 2940.450 839.730 2943.350 839.790 ;
        RECT -23.730 836.830 2943.350 839.730 ;
        RECT -23.730 836.770 -20.830 836.830 ;
        RECT 111.470 836.770 114.370 836.830 ;
        RECT 291.470 836.770 294.370 836.830 ;
        RECT 471.470 836.770 474.370 836.830 ;
        RECT 651.470 836.770 654.370 836.830 ;
        RECT 831.470 836.770 834.370 836.830 ;
        RECT 1011.470 836.770 1014.370 836.830 ;
        RECT 1191.470 836.770 1194.370 836.830 ;
        RECT 1371.470 836.770 1374.370 836.830 ;
        RECT 1551.470 836.770 1554.370 836.830 ;
        RECT 1731.470 836.770 1734.370 836.830 ;
        RECT 1911.470 836.770 1914.370 836.830 ;
        RECT 2091.470 836.770 2094.370 836.830 ;
        RECT 2271.470 836.770 2274.370 836.830 ;
        RECT 2451.470 836.770 2454.370 836.830 ;
        RECT 2631.470 836.770 2634.370 836.830 ;
        RECT 2811.470 836.770 2814.370 836.830 ;
        RECT 2940.450 836.770 2943.350 836.830 ;
        RECT -23.730 659.730 -20.830 659.790 ;
        RECT 111.470 659.730 114.370 659.790 ;
        RECT 291.470 659.730 294.370 659.790 ;
        RECT 471.470 659.730 474.370 659.790 ;
        RECT 651.470 659.730 654.370 659.790 ;
        RECT 831.470 659.730 834.370 659.790 ;
        RECT 1011.470 659.730 1014.370 659.790 ;
        RECT 1191.470 659.730 1194.370 659.790 ;
        RECT 1371.470 659.730 1374.370 659.790 ;
        RECT 1551.470 659.730 1554.370 659.790 ;
        RECT 1731.470 659.730 1734.370 659.790 ;
        RECT 1911.470 659.730 1914.370 659.790 ;
        RECT 2091.470 659.730 2094.370 659.790 ;
        RECT 2271.470 659.730 2274.370 659.790 ;
        RECT 2451.470 659.730 2454.370 659.790 ;
        RECT 2631.470 659.730 2634.370 659.790 ;
        RECT 2811.470 659.730 2814.370 659.790 ;
        RECT 2940.450 659.730 2943.350 659.790 ;
        RECT -23.730 656.830 2943.350 659.730 ;
        RECT -23.730 656.770 -20.830 656.830 ;
        RECT 111.470 656.770 114.370 656.830 ;
        RECT 291.470 656.770 294.370 656.830 ;
        RECT 471.470 656.770 474.370 656.830 ;
        RECT 651.470 656.770 654.370 656.830 ;
        RECT 831.470 656.770 834.370 656.830 ;
        RECT 1011.470 656.770 1014.370 656.830 ;
        RECT 1191.470 656.770 1194.370 656.830 ;
        RECT 1371.470 656.770 1374.370 656.830 ;
        RECT 1551.470 656.770 1554.370 656.830 ;
        RECT 1731.470 656.770 1734.370 656.830 ;
        RECT 1911.470 656.770 1914.370 656.830 ;
        RECT 2091.470 656.770 2094.370 656.830 ;
        RECT 2271.470 656.770 2274.370 656.830 ;
        RECT 2451.470 656.770 2454.370 656.830 ;
        RECT 2631.470 656.770 2634.370 656.830 ;
        RECT 2811.470 656.770 2814.370 656.830 ;
        RECT 2940.450 656.770 2943.350 656.830 ;
        RECT -23.730 479.730 -20.830 479.790 ;
        RECT 111.470 479.730 114.370 479.790 ;
        RECT 291.470 479.730 294.370 479.790 ;
        RECT 471.470 479.730 474.370 479.790 ;
        RECT 651.470 479.730 654.370 479.790 ;
        RECT 831.470 479.730 834.370 479.790 ;
        RECT 1011.470 479.730 1014.370 479.790 ;
        RECT 1191.470 479.730 1194.370 479.790 ;
        RECT 1371.470 479.730 1374.370 479.790 ;
        RECT 1551.470 479.730 1554.370 479.790 ;
        RECT 1731.470 479.730 1734.370 479.790 ;
        RECT 1911.470 479.730 1914.370 479.790 ;
        RECT 2091.470 479.730 2094.370 479.790 ;
        RECT 2271.470 479.730 2274.370 479.790 ;
        RECT 2451.470 479.730 2454.370 479.790 ;
        RECT 2631.470 479.730 2634.370 479.790 ;
        RECT 2811.470 479.730 2814.370 479.790 ;
        RECT 2940.450 479.730 2943.350 479.790 ;
        RECT -23.730 476.830 2943.350 479.730 ;
        RECT -23.730 476.770 -20.830 476.830 ;
        RECT 111.470 476.770 114.370 476.830 ;
        RECT 291.470 476.770 294.370 476.830 ;
        RECT 471.470 476.770 474.370 476.830 ;
        RECT 651.470 476.770 654.370 476.830 ;
        RECT 831.470 476.770 834.370 476.830 ;
        RECT 1011.470 476.770 1014.370 476.830 ;
        RECT 1191.470 476.770 1194.370 476.830 ;
        RECT 1371.470 476.770 1374.370 476.830 ;
        RECT 1551.470 476.770 1554.370 476.830 ;
        RECT 1731.470 476.770 1734.370 476.830 ;
        RECT 1911.470 476.770 1914.370 476.830 ;
        RECT 2091.470 476.770 2094.370 476.830 ;
        RECT 2271.470 476.770 2274.370 476.830 ;
        RECT 2451.470 476.770 2454.370 476.830 ;
        RECT 2631.470 476.770 2634.370 476.830 ;
        RECT 2811.470 476.770 2814.370 476.830 ;
        RECT 2940.450 476.770 2943.350 476.830 ;
        RECT -23.730 299.730 -20.830 299.790 ;
        RECT 111.470 299.730 114.370 299.790 ;
        RECT 291.470 299.730 294.370 299.790 ;
        RECT 471.470 299.730 474.370 299.790 ;
        RECT 651.470 299.730 654.370 299.790 ;
        RECT 831.470 299.730 834.370 299.790 ;
        RECT 1011.470 299.730 1014.370 299.790 ;
        RECT 1191.470 299.730 1194.370 299.790 ;
        RECT 1371.470 299.730 1374.370 299.790 ;
        RECT 1551.470 299.730 1554.370 299.790 ;
        RECT 1731.470 299.730 1734.370 299.790 ;
        RECT 1911.470 299.730 1914.370 299.790 ;
        RECT 2091.470 299.730 2094.370 299.790 ;
        RECT 2271.470 299.730 2274.370 299.790 ;
        RECT 2451.470 299.730 2454.370 299.790 ;
        RECT 2631.470 299.730 2634.370 299.790 ;
        RECT 2811.470 299.730 2814.370 299.790 ;
        RECT 2940.450 299.730 2943.350 299.790 ;
        RECT -23.730 296.830 2943.350 299.730 ;
        RECT -23.730 296.770 -20.830 296.830 ;
        RECT 111.470 296.770 114.370 296.830 ;
        RECT 291.470 296.770 294.370 296.830 ;
        RECT 471.470 296.770 474.370 296.830 ;
        RECT 651.470 296.770 654.370 296.830 ;
        RECT 831.470 296.770 834.370 296.830 ;
        RECT 1011.470 296.770 1014.370 296.830 ;
        RECT 1191.470 296.770 1194.370 296.830 ;
        RECT 1371.470 296.770 1374.370 296.830 ;
        RECT 1551.470 296.770 1554.370 296.830 ;
        RECT 1731.470 296.770 1734.370 296.830 ;
        RECT 1911.470 296.770 1914.370 296.830 ;
        RECT 2091.470 296.770 2094.370 296.830 ;
        RECT 2271.470 296.770 2274.370 296.830 ;
        RECT 2451.470 296.770 2454.370 296.830 ;
        RECT 2631.470 296.770 2634.370 296.830 ;
        RECT 2811.470 296.770 2814.370 296.830 ;
        RECT 2940.450 296.770 2943.350 296.830 ;
        RECT -23.730 119.730 -20.830 119.790 ;
        RECT 111.470 119.730 114.370 119.790 ;
        RECT 291.470 119.730 294.370 119.790 ;
        RECT 471.470 119.730 474.370 119.790 ;
        RECT 651.470 119.730 654.370 119.790 ;
        RECT 831.470 119.730 834.370 119.790 ;
        RECT 1011.470 119.730 1014.370 119.790 ;
        RECT 1191.470 119.730 1194.370 119.790 ;
        RECT 1371.470 119.730 1374.370 119.790 ;
        RECT 1551.470 119.730 1554.370 119.790 ;
        RECT 1731.470 119.730 1734.370 119.790 ;
        RECT 1911.470 119.730 1914.370 119.790 ;
        RECT 2091.470 119.730 2094.370 119.790 ;
        RECT 2271.470 119.730 2274.370 119.790 ;
        RECT 2451.470 119.730 2454.370 119.790 ;
        RECT 2631.470 119.730 2634.370 119.790 ;
        RECT 2811.470 119.730 2814.370 119.790 ;
        RECT 2940.450 119.730 2943.350 119.790 ;
        RECT -23.730 116.830 2943.350 119.730 ;
        RECT -23.730 116.770 -20.830 116.830 ;
        RECT 111.470 116.770 114.370 116.830 ;
        RECT 291.470 116.770 294.370 116.830 ;
        RECT 471.470 116.770 474.370 116.830 ;
        RECT 651.470 116.770 654.370 116.830 ;
        RECT 831.470 116.770 834.370 116.830 ;
        RECT 1011.470 116.770 1014.370 116.830 ;
        RECT 1191.470 116.770 1194.370 116.830 ;
        RECT 1371.470 116.770 1374.370 116.830 ;
        RECT 1551.470 116.770 1554.370 116.830 ;
        RECT 1731.470 116.770 1734.370 116.830 ;
        RECT 1911.470 116.770 1914.370 116.830 ;
        RECT 2091.470 116.770 2094.370 116.830 ;
        RECT 2271.470 116.770 2274.370 116.830 ;
        RECT 2451.470 116.770 2454.370 116.830 ;
        RECT 2631.470 116.770 2634.370 116.830 ;
        RECT 2811.470 116.770 2814.370 116.830 ;
        RECT 2940.450 116.770 2943.350 116.830 ;
        RECT -23.730 -15.470 -20.830 -15.410 ;
        RECT 111.470 -15.470 114.370 -15.410 ;
        RECT 291.470 -15.470 294.370 -15.410 ;
        RECT 471.470 -15.470 474.370 -15.410 ;
        RECT 651.470 -15.470 654.370 -15.410 ;
        RECT 831.470 -15.470 834.370 -15.410 ;
        RECT 1011.470 -15.470 1014.370 -15.410 ;
        RECT 1191.470 -15.470 1194.370 -15.410 ;
        RECT 1371.470 -15.470 1374.370 -15.410 ;
        RECT 1551.470 -15.470 1554.370 -15.410 ;
        RECT 1731.470 -15.470 1734.370 -15.410 ;
        RECT 1911.470 -15.470 1914.370 -15.410 ;
        RECT 2091.470 -15.470 2094.370 -15.410 ;
        RECT 2271.470 -15.470 2274.370 -15.410 ;
        RECT 2451.470 -15.470 2454.370 -15.410 ;
        RECT 2631.470 -15.470 2634.370 -15.410 ;
        RECT 2811.470 -15.470 2814.370 -15.410 ;
        RECT 2940.450 -15.470 2943.350 -15.410 ;
        RECT -23.730 -18.370 2943.350 -15.470 ;
        RECT -23.730 -18.430 -20.830 -18.370 ;
        RECT 111.470 -18.430 114.370 -18.370 ;
        RECT 291.470 -18.430 294.370 -18.370 ;
        RECT 471.470 -18.430 474.370 -18.370 ;
        RECT 651.470 -18.430 654.370 -18.370 ;
        RECT 831.470 -18.430 834.370 -18.370 ;
        RECT 1011.470 -18.430 1014.370 -18.370 ;
        RECT 1191.470 -18.430 1194.370 -18.370 ;
        RECT 1371.470 -18.430 1374.370 -18.370 ;
        RECT 1551.470 -18.430 1554.370 -18.370 ;
        RECT 1731.470 -18.430 1734.370 -18.370 ;
        RECT 1911.470 -18.430 1914.370 -18.370 ;
        RECT 2091.470 -18.430 2094.370 -18.370 ;
        RECT 2271.470 -18.430 2274.370 -18.370 ;
        RECT 2451.470 -18.430 2454.370 -18.370 ;
        RECT 2631.470 -18.430 2634.370 -18.370 ;
        RECT 2811.470 -18.430 2814.370 -18.370 ;
        RECT 2940.450 -18.430 2943.350 -18.370 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.330 -22.970 -25.430 3542.650 ;
        RECT 38.870 -27.570 41.770 3547.250 ;
        RECT 218.870 -27.570 221.770 3547.250 ;
        RECT 398.870 -27.570 401.770 3547.250 ;
        RECT 578.870 -27.570 581.770 3547.250 ;
        RECT 758.870 -27.570 761.770 3547.250 ;
        RECT 938.870 -27.570 941.770 3547.250 ;
        RECT 1118.870 -27.570 1121.770 3547.250 ;
        RECT 1298.870 -27.570 1301.770 3547.250 ;
        RECT 1478.870 -27.570 1481.770 3547.250 ;
        RECT 1658.870 -27.570 1661.770 3547.250 ;
        RECT 1838.870 -27.570 1841.770 3547.250 ;
        RECT 2018.870 -27.570 2021.770 3547.250 ;
        RECT 2198.870 -27.570 2201.770 3547.250 ;
        RECT 2378.870 -27.570 2381.770 3547.250 ;
        RECT 2558.870 -27.570 2561.770 3547.250 ;
        RECT 2738.870 -27.570 2741.770 3547.250 ;
        RECT 2945.050 -22.970 2947.950 3542.650 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3465.890 -26.290 3467.070 ;
        RECT -27.470 3464.290 -26.290 3465.470 ;
        RECT -27.470 3285.890 -26.290 3287.070 ;
        RECT -27.470 3284.290 -26.290 3285.470 ;
        RECT -27.470 3105.890 -26.290 3107.070 ;
        RECT -27.470 3104.290 -26.290 3105.470 ;
        RECT -27.470 2925.890 -26.290 2927.070 ;
        RECT -27.470 2924.290 -26.290 2925.470 ;
        RECT -27.470 2745.890 -26.290 2747.070 ;
        RECT -27.470 2744.290 -26.290 2745.470 ;
        RECT -27.470 2565.890 -26.290 2567.070 ;
        RECT -27.470 2564.290 -26.290 2565.470 ;
        RECT -27.470 2385.890 -26.290 2387.070 ;
        RECT -27.470 2384.290 -26.290 2385.470 ;
        RECT -27.470 2205.890 -26.290 2207.070 ;
        RECT -27.470 2204.290 -26.290 2205.470 ;
        RECT -27.470 2025.890 -26.290 2027.070 ;
        RECT -27.470 2024.290 -26.290 2025.470 ;
        RECT -27.470 1845.890 -26.290 1847.070 ;
        RECT -27.470 1844.290 -26.290 1845.470 ;
        RECT -27.470 1665.890 -26.290 1667.070 ;
        RECT -27.470 1664.290 -26.290 1665.470 ;
        RECT -27.470 1485.890 -26.290 1487.070 ;
        RECT -27.470 1484.290 -26.290 1485.470 ;
        RECT -27.470 1305.890 -26.290 1307.070 ;
        RECT -27.470 1304.290 -26.290 1305.470 ;
        RECT -27.470 1125.890 -26.290 1127.070 ;
        RECT -27.470 1124.290 -26.290 1125.470 ;
        RECT -27.470 945.890 -26.290 947.070 ;
        RECT -27.470 944.290 -26.290 945.470 ;
        RECT -27.470 765.890 -26.290 767.070 ;
        RECT -27.470 764.290 -26.290 765.470 ;
        RECT -27.470 585.890 -26.290 587.070 ;
        RECT -27.470 584.290 -26.290 585.470 ;
        RECT -27.470 405.890 -26.290 407.070 ;
        RECT -27.470 404.290 -26.290 405.470 ;
        RECT -27.470 225.890 -26.290 227.070 ;
        RECT -27.470 224.290 -26.290 225.470 ;
        RECT -27.470 45.890 -26.290 47.070 ;
        RECT -27.470 44.290 -26.290 45.470 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 39.730 3541.410 40.910 3542.590 ;
        RECT 39.730 3539.810 40.910 3540.990 ;
        RECT 39.730 3465.890 40.910 3467.070 ;
        RECT 39.730 3464.290 40.910 3465.470 ;
        RECT 39.730 3285.890 40.910 3287.070 ;
        RECT 39.730 3284.290 40.910 3285.470 ;
        RECT 39.730 3105.890 40.910 3107.070 ;
        RECT 39.730 3104.290 40.910 3105.470 ;
        RECT 39.730 2925.890 40.910 2927.070 ;
        RECT 39.730 2924.290 40.910 2925.470 ;
        RECT 39.730 2745.890 40.910 2747.070 ;
        RECT 39.730 2744.290 40.910 2745.470 ;
        RECT 39.730 2565.890 40.910 2567.070 ;
        RECT 39.730 2564.290 40.910 2565.470 ;
        RECT 39.730 2385.890 40.910 2387.070 ;
        RECT 39.730 2384.290 40.910 2385.470 ;
        RECT 39.730 2205.890 40.910 2207.070 ;
        RECT 39.730 2204.290 40.910 2205.470 ;
        RECT 39.730 2025.890 40.910 2027.070 ;
        RECT 39.730 2024.290 40.910 2025.470 ;
        RECT 39.730 1845.890 40.910 1847.070 ;
        RECT 39.730 1844.290 40.910 1845.470 ;
        RECT 39.730 1665.890 40.910 1667.070 ;
        RECT 39.730 1664.290 40.910 1665.470 ;
        RECT 39.730 1485.890 40.910 1487.070 ;
        RECT 39.730 1484.290 40.910 1485.470 ;
        RECT 39.730 1305.890 40.910 1307.070 ;
        RECT 39.730 1304.290 40.910 1305.470 ;
        RECT 39.730 1125.890 40.910 1127.070 ;
        RECT 39.730 1124.290 40.910 1125.470 ;
        RECT 39.730 945.890 40.910 947.070 ;
        RECT 39.730 944.290 40.910 945.470 ;
        RECT 39.730 765.890 40.910 767.070 ;
        RECT 39.730 764.290 40.910 765.470 ;
        RECT 39.730 585.890 40.910 587.070 ;
        RECT 39.730 584.290 40.910 585.470 ;
        RECT 39.730 405.890 40.910 407.070 ;
        RECT 39.730 404.290 40.910 405.470 ;
        RECT 39.730 225.890 40.910 227.070 ;
        RECT 39.730 224.290 40.910 225.470 ;
        RECT 39.730 45.890 40.910 47.070 ;
        RECT 39.730 44.290 40.910 45.470 ;
        RECT 39.730 -21.310 40.910 -20.130 ;
        RECT 39.730 -22.910 40.910 -21.730 ;
        RECT 219.730 3541.410 220.910 3542.590 ;
        RECT 219.730 3539.810 220.910 3540.990 ;
        RECT 219.730 3465.890 220.910 3467.070 ;
        RECT 219.730 3464.290 220.910 3465.470 ;
        RECT 219.730 3285.890 220.910 3287.070 ;
        RECT 219.730 3284.290 220.910 3285.470 ;
        RECT 219.730 3105.890 220.910 3107.070 ;
        RECT 219.730 3104.290 220.910 3105.470 ;
        RECT 219.730 2925.890 220.910 2927.070 ;
        RECT 219.730 2924.290 220.910 2925.470 ;
        RECT 219.730 2745.890 220.910 2747.070 ;
        RECT 219.730 2744.290 220.910 2745.470 ;
        RECT 219.730 2565.890 220.910 2567.070 ;
        RECT 219.730 2564.290 220.910 2565.470 ;
        RECT 219.730 2385.890 220.910 2387.070 ;
        RECT 219.730 2384.290 220.910 2385.470 ;
        RECT 219.730 2205.890 220.910 2207.070 ;
        RECT 219.730 2204.290 220.910 2205.470 ;
        RECT 219.730 2025.890 220.910 2027.070 ;
        RECT 219.730 2024.290 220.910 2025.470 ;
        RECT 219.730 1845.890 220.910 1847.070 ;
        RECT 219.730 1844.290 220.910 1845.470 ;
        RECT 219.730 1665.890 220.910 1667.070 ;
        RECT 219.730 1664.290 220.910 1665.470 ;
        RECT 219.730 1485.890 220.910 1487.070 ;
        RECT 219.730 1484.290 220.910 1485.470 ;
        RECT 219.730 1305.890 220.910 1307.070 ;
        RECT 219.730 1304.290 220.910 1305.470 ;
        RECT 219.730 1125.890 220.910 1127.070 ;
        RECT 219.730 1124.290 220.910 1125.470 ;
        RECT 219.730 945.890 220.910 947.070 ;
        RECT 219.730 944.290 220.910 945.470 ;
        RECT 219.730 765.890 220.910 767.070 ;
        RECT 219.730 764.290 220.910 765.470 ;
        RECT 219.730 585.890 220.910 587.070 ;
        RECT 219.730 584.290 220.910 585.470 ;
        RECT 219.730 405.890 220.910 407.070 ;
        RECT 219.730 404.290 220.910 405.470 ;
        RECT 219.730 225.890 220.910 227.070 ;
        RECT 219.730 224.290 220.910 225.470 ;
        RECT 219.730 45.890 220.910 47.070 ;
        RECT 219.730 44.290 220.910 45.470 ;
        RECT 219.730 -21.310 220.910 -20.130 ;
        RECT 219.730 -22.910 220.910 -21.730 ;
        RECT 399.730 3541.410 400.910 3542.590 ;
        RECT 399.730 3539.810 400.910 3540.990 ;
        RECT 399.730 3465.890 400.910 3467.070 ;
        RECT 399.730 3464.290 400.910 3465.470 ;
        RECT 399.730 3285.890 400.910 3287.070 ;
        RECT 399.730 3284.290 400.910 3285.470 ;
        RECT 399.730 3105.890 400.910 3107.070 ;
        RECT 399.730 3104.290 400.910 3105.470 ;
        RECT 399.730 2925.890 400.910 2927.070 ;
        RECT 399.730 2924.290 400.910 2925.470 ;
        RECT 399.730 2745.890 400.910 2747.070 ;
        RECT 399.730 2744.290 400.910 2745.470 ;
        RECT 399.730 2565.890 400.910 2567.070 ;
        RECT 399.730 2564.290 400.910 2565.470 ;
        RECT 399.730 2385.890 400.910 2387.070 ;
        RECT 399.730 2384.290 400.910 2385.470 ;
        RECT 399.730 2205.890 400.910 2207.070 ;
        RECT 399.730 2204.290 400.910 2205.470 ;
        RECT 399.730 2025.890 400.910 2027.070 ;
        RECT 399.730 2024.290 400.910 2025.470 ;
        RECT 399.730 1845.890 400.910 1847.070 ;
        RECT 399.730 1844.290 400.910 1845.470 ;
        RECT 399.730 1665.890 400.910 1667.070 ;
        RECT 399.730 1664.290 400.910 1665.470 ;
        RECT 399.730 1485.890 400.910 1487.070 ;
        RECT 399.730 1484.290 400.910 1485.470 ;
        RECT 399.730 1305.890 400.910 1307.070 ;
        RECT 399.730 1304.290 400.910 1305.470 ;
        RECT 399.730 1125.890 400.910 1127.070 ;
        RECT 399.730 1124.290 400.910 1125.470 ;
        RECT 399.730 945.890 400.910 947.070 ;
        RECT 399.730 944.290 400.910 945.470 ;
        RECT 399.730 765.890 400.910 767.070 ;
        RECT 399.730 764.290 400.910 765.470 ;
        RECT 399.730 585.890 400.910 587.070 ;
        RECT 399.730 584.290 400.910 585.470 ;
        RECT 399.730 405.890 400.910 407.070 ;
        RECT 399.730 404.290 400.910 405.470 ;
        RECT 399.730 225.890 400.910 227.070 ;
        RECT 399.730 224.290 400.910 225.470 ;
        RECT 399.730 45.890 400.910 47.070 ;
        RECT 399.730 44.290 400.910 45.470 ;
        RECT 399.730 -21.310 400.910 -20.130 ;
        RECT 399.730 -22.910 400.910 -21.730 ;
        RECT 579.730 3541.410 580.910 3542.590 ;
        RECT 579.730 3539.810 580.910 3540.990 ;
        RECT 579.730 3465.890 580.910 3467.070 ;
        RECT 579.730 3464.290 580.910 3465.470 ;
        RECT 579.730 3285.890 580.910 3287.070 ;
        RECT 579.730 3284.290 580.910 3285.470 ;
        RECT 579.730 3105.890 580.910 3107.070 ;
        RECT 579.730 3104.290 580.910 3105.470 ;
        RECT 579.730 2925.890 580.910 2927.070 ;
        RECT 579.730 2924.290 580.910 2925.470 ;
        RECT 579.730 2745.890 580.910 2747.070 ;
        RECT 579.730 2744.290 580.910 2745.470 ;
        RECT 579.730 2565.890 580.910 2567.070 ;
        RECT 579.730 2564.290 580.910 2565.470 ;
        RECT 579.730 2385.890 580.910 2387.070 ;
        RECT 579.730 2384.290 580.910 2385.470 ;
        RECT 579.730 2205.890 580.910 2207.070 ;
        RECT 579.730 2204.290 580.910 2205.470 ;
        RECT 579.730 2025.890 580.910 2027.070 ;
        RECT 579.730 2024.290 580.910 2025.470 ;
        RECT 579.730 1845.890 580.910 1847.070 ;
        RECT 579.730 1844.290 580.910 1845.470 ;
        RECT 579.730 1665.890 580.910 1667.070 ;
        RECT 579.730 1664.290 580.910 1665.470 ;
        RECT 579.730 1485.890 580.910 1487.070 ;
        RECT 579.730 1484.290 580.910 1485.470 ;
        RECT 579.730 1305.890 580.910 1307.070 ;
        RECT 579.730 1304.290 580.910 1305.470 ;
        RECT 579.730 1125.890 580.910 1127.070 ;
        RECT 579.730 1124.290 580.910 1125.470 ;
        RECT 579.730 945.890 580.910 947.070 ;
        RECT 579.730 944.290 580.910 945.470 ;
        RECT 579.730 765.890 580.910 767.070 ;
        RECT 579.730 764.290 580.910 765.470 ;
        RECT 579.730 585.890 580.910 587.070 ;
        RECT 579.730 584.290 580.910 585.470 ;
        RECT 579.730 405.890 580.910 407.070 ;
        RECT 579.730 404.290 580.910 405.470 ;
        RECT 579.730 225.890 580.910 227.070 ;
        RECT 579.730 224.290 580.910 225.470 ;
        RECT 579.730 45.890 580.910 47.070 ;
        RECT 579.730 44.290 580.910 45.470 ;
        RECT 579.730 -21.310 580.910 -20.130 ;
        RECT 579.730 -22.910 580.910 -21.730 ;
        RECT 759.730 3541.410 760.910 3542.590 ;
        RECT 759.730 3539.810 760.910 3540.990 ;
        RECT 759.730 3465.890 760.910 3467.070 ;
        RECT 759.730 3464.290 760.910 3465.470 ;
        RECT 759.730 3285.890 760.910 3287.070 ;
        RECT 759.730 3284.290 760.910 3285.470 ;
        RECT 759.730 3105.890 760.910 3107.070 ;
        RECT 759.730 3104.290 760.910 3105.470 ;
        RECT 759.730 2925.890 760.910 2927.070 ;
        RECT 759.730 2924.290 760.910 2925.470 ;
        RECT 759.730 2745.890 760.910 2747.070 ;
        RECT 759.730 2744.290 760.910 2745.470 ;
        RECT 759.730 2565.890 760.910 2567.070 ;
        RECT 759.730 2564.290 760.910 2565.470 ;
        RECT 759.730 2385.890 760.910 2387.070 ;
        RECT 759.730 2384.290 760.910 2385.470 ;
        RECT 759.730 2205.890 760.910 2207.070 ;
        RECT 759.730 2204.290 760.910 2205.470 ;
        RECT 759.730 2025.890 760.910 2027.070 ;
        RECT 759.730 2024.290 760.910 2025.470 ;
        RECT 759.730 1845.890 760.910 1847.070 ;
        RECT 759.730 1844.290 760.910 1845.470 ;
        RECT 759.730 1665.890 760.910 1667.070 ;
        RECT 759.730 1664.290 760.910 1665.470 ;
        RECT 759.730 1485.890 760.910 1487.070 ;
        RECT 759.730 1484.290 760.910 1485.470 ;
        RECT 759.730 1305.890 760.910 1307.070 ;
        RECT 759.730 1304.290 760.910 1305.470 ;
        RECT 759.730 1125.890 760.910 1127.070 ;
        RECT 759.730 1124.290 760.910 1125.470 ;
        RECT 759.730 945.890 760.910 947.070 ;
        RECT 759.730 944.290 760.910 945.470 ;
        RECT 759.730 765.890 760.910 767.070 ;
        RECT 759.730 764.290 760.910 765.470 ;
        RECT 759.730 585.890 760.910 587.070 ;
        RECT 759.730 584.290 760.910 585.470 ;
        RECT 759.730 405.890 760.910 407.070 ;
        RECT 759.730 404.290 760.910 405.470 ;
        RECT 759.730 225.890 760.910 227.070 ;
        RECT 759.730 224.290 760.910 225.470 ;
        RECT 759.730 45.890 760.910 47.070 ;
        RECT 759.730 44.290 760.910 45.470 ;
        RECT 759.730 -21.310 760.910 -20.130 ;
        RECT 759.730 -22.910 760.910 -21.730 ;
        RECT 939.730 3541.410 940.910 3542.590 ;
        RECT 939.730 3539.810 940.910 3540.990 ;
        RECT 939.730 3465.890 940.910 3467.070 ;
        RECT 939.730 3464.290 940.910 3465.470 ;
        RECT 939.730 3285.890 940.910 3287.070 ;
        RECT 939.730 3284.290 940.910 3285.470 ;
        RECT 939.730 3105.890 940.910 3107.070 ;
        RECT 939.730 3104.290 940.910 3105.470 ;
        RECT 939.730 2925.890 940.910 2927.070 ;
        RECT 939.730 2924.290 940.910 2925.470 ;
        RECT 939.730 2745.890 940.910 2747.070 ;
        RECT 939.730 2744.290 940.910 2745.470 ;
        RECT 939.730 2565.890 940.910 2567.070 ;
        RECT 939.730 2564.290 940.910 2565.470 ;
        RECT 939.730 2385.890 940.910 2387.070 ;
        RECT 939.730 2384.290 940.910 2385.470 ;
        RECT 939.730 2205.890 940.910 2207.070 ;
        RECT 939.730 2204.290 940.910 2205.470 ;
        RECT 939.730 2025.890 940.910 2027.070 ;
        RECT 939.730 2024.290 940.910 2025.470 ;
        RECT 939.730 1845.890 940.910 1847.070 ;
        RECT 939.730 1844.290 940.910 1845.470 ;
        RECT 939.730 1665.890 940.910 1667.070 ;
        RECT 939.730 1664.290 940.910 1665.470 ;
        RECT 939.730 1485.890 940.910 1487.070 ;
        RECT 939.730 1484.290 940.910 1485.470 ;
        RECT 939.730 1305.890 940.910 1307.070 ;
        RECT 939.730 1304.290 940.910 1305.470 ;
        RECT 939.730 1125.890 940.910 1127.070 ;
        RECT 939.730 1124.290 940.910 1125.470 ;
        RECT 939.730 945.890 940.910 947.070 ;
        RECT 939.730 944.290 940.910 945.470 ;
        RECT 939.730 765.890 940.910 767.070 ;
        RECT 939.730 764.290 940.910 765.470 ;
        RECT 939.730 585.890 940.910 587.070 ;
        RECT 939.730 584.290 940.910 585.470 ;
        RECT 939.730 405.890 940.910 407.070 ;
        RECT 939.730 404.290 940.910 405.470 ;
        RECT 939.730 225.890 940.910 227.070 ;
        RECT 939.730 224.290 940.910 225.470 ;
        RECT 939.730 45.890 940.910 47.070 ;
        RECT 939.730 44.290 940.910 45.470 ;
        RECT 939.730 -21.310 940.910 -20.130 ;
        RECT 939.730 -22.910 940.910 -21.730 ;
        RECT 1119.730 3541.410 1120.910 3542.590 ;
        RECT 1119.730 3539.810 1120.910 3540.990 ;
        RECT 1119.730 3465.890 1120.910 3467.070 ;
        RECT 1119.730 3464.290 1120.910 3465.470 ;
        RECT 1119.730 3285.890 1120.910 3287.070 ;
        RECT 1119.730 3284.290 1120.910 3285.470 ;
        RECT 1119.730 3105.890 1120.910 3107.070 ;
        RECT 1119.730 3104.290 1120.910 3105.470 ;
        RECT 1119.730 2925.890 1120.910 2927.070 ;
        RECT 1119.730 2924.290 1120.910 2925.470 ;
        RECT 1119.730 2745.890 1120.910 2747.070 ;
        RECT 1119.730 2744.290 1120.910 2745.470 ;
        RECT 1119.730 2565.890 1120.910 2567.070 ;
        RECT 1119.730 2564.290 1120.910 2565.470 ;
        RECT 1119.730 2385.890 1120.910 2387.070 ;
        RECT 1119.730 2384.290 1120.910 2385.470 ;
        RECT 1119.730 2205.890 1120.910 2207.070 ;
        RECT 1119.730 2204.290 1120.910 2205.470 ;
        RECT 1119.730 2025.890 1120.910 2027.070 ;
        RECT 1119.730 2024.290 1120.910 2025.470 ;
        RECT 1119.730 1845.890 1120.910 1847.070 ;
        RECT 1119.730 1844.290 1120.910 1845.470 ;
        RECT 1119.730 1665.890 1120.910 1667.070 ;
        RECT 1119.730 1664.290 1120.910 1665.470 ;
        RECT 1119.730 1485.890 1120.910 1487.070 ;
        RECT 1119.730 1484.290 1120.910 1485.470 ;
        RECT 1119.730 1305.890 1120.910 1307.070 ;
        RECT 1119.730 1304.290 1120.910 1305.470 ;
        RECT 1119.730 1125.890 1120.910 1127.070 ;
        RECT 1119.730 1124.290 1120.910 1125.470 ;
        RECT 1119.730 945.890 1120.910 947.070 ;
        RECT 1119.730 944.290 1120.910 945.470 ;
        RECT 1119.730 765.890 1120.910 767.070 ;
        RECT 1119.730 764.290 1120.910 765.470 ;
        RECT 1119.730 585.890 1120.910 587.070 ;
        RECT 1119.730 584.290 1120.910 585.470 ;
        RECT 1119.730 405.890 1120.910 407.070 ;
        RECT 1119.730 404.290 1120.910 405.470 ;
        RECT 1119.730 225.890 1120.910 227.070 ;
        RECT 1119.730 224.290 1120.910 225.470 ;
        RECT 1119.730 45.890 1120.910 47.070 ;
        RECT 1119.730 44.290 1120.910 45.470 ;
        RECT 1119.730 -21.310 1120.910 -20.130 ;
        RECT 1119.730 -22.910 1120.910 -21.730 ;
        RECT 1299.730 3541.410 1300.910 3542.590 ;
        RECT 1299.730 3539.810 1300.910 3540.990 ;
        RECT 1299.730 3465.890 1300.910 3467.070 ;
        RECT 1299.730 3464.290 1300.910 3465.470 ;
        RECT 1299.730 3285.890 1300.910 3287.070 ;
        RECT 1299.730 3284.290 1300.910 3285.470 ;
        RECT 1299.730 3105.890 1300.910 3107.070 ;
        RECT 1299.730 3104.290 1300.910 3105.470 ;
        RECT 1299.730 2925.890 1300.910 2927.070 ;
        RECT 1299.730 2924.290 1300.910 2925.470 ;
        RECT 1299.730 2745.890 1300.910 2747.070 ;
        RECT 1299.730 2744.290 1300.910 2745.470 ;
        RECT 1299.730 2565.890 1300.910 2567.070 ;
        RECT 1299.730 2564.290 1300.910 2565.470 ;
        RECT 1299.730 2385.890 1300.910 2387.070 ;
        RECT 1299.730 2384.290 1300.910 2385.470 ;
        RECT 1299.730 2205.890 1300.910 2207.070 ;
        RECT 1299.730 2204.290 1300.910 2205.470 ;
        RECT 1299.730 2025.890 1300.910 2027.070 ;
        RECT 1299.730 2024.290 1300.910 2025.470 ;
        RECT 1299.730 1845.890 1300.910 1847.070 ;
        RECT 1299.730 1844.290 1300.910 1845.470 ;
        RECT 1299.730 1665.890 1300.910 1667.070 ;
        RECT 1299.730 1664.290 1300.910 1665.470 ;
        RECT 1299.730 1485.890 1300.910 1487.070 ;
        RECT 1299.730 1484.290 1300.910 1485.470 ;
        RECT 1299.730 1305.890 1300.910 1307.070 ;
        RECT 1299.730 1304.290 1300.910 1305.470 ;
        RECT 1299.730 1125.890 1300.910 1127.070 ;
        RECT 1299.730 1124.290 1300.910 1125.470 ;
        RECT 1299.730 945.890 1300.910 947.070 ;
        RECT 1299.730 944.290 1300.910 945.470 ;
        RECT 1299.730 765.890 1300.910 767.070 ;
        RECT 1299.730 764.290 1300.910 765.470 ;
        RECT 1299.730 585.890 1300.910 587.070 ;
        RECT 1299.730 584.290 1300.910 585.470 ;
        RECT 1299.730 405.890 1300.910 407.070 ;
        RECT 1299.730 404.290 1300.910 405.470 ;
        RECT 1299.730 225.890 1300.910 227.070 ;
        RECT 1299.730 224.290 1300.910 225.470 ;
        RECT 1299.730 45.890 1300.910 47.070 ;
        RECT 1299.730 44.290 1300.910 45.470 ;
        RECT 1299.730 -21.310 1300.910 -20.130 ;
        RECT 1299.730 -22.910 1300.910 -21.730 ;
        RECT 1479.730 3541.410 1480.910 3542.590 ;
        RECT 1479.730 3539.810 1480.910 3540.990 ;
        RECT 1479.730 3465.890 1480.910 3467.070 ;
        RECT 1479.730 3464.290 1480.910 3465.470 ;
        RECT 1479.730 3285.890 1480.910 3287.070 ;
        RECT 1479.730 3284.290 1480.910 3285.470 ;
        RECT 1479.730 3105.890 1480.910 3107.070 ;
        RECT 1479.730 3104.290 1480.910 3105.470 ;
        RECT 1479.730 2925.890 1480.910 2927.070 ;
        RECT 1479.730 2924.290 1480.910 2925.470 ;
        RECT 1479.730 2745.890 1480.910 2747.070 ;
        RECT 1479.730 2744.290 1480.910 2745.470 ;
        RECT 1479.730 2565.890 1480.910 2567.070 ;
        RECT 1479.730 2564.290 1480.910 2565.470 ;
        RECT 1479.730 2385.890 1480.910 2387.070 ;
        RECT 1479.730 2384.290 1480.910 2385.470 ;
        RECT 1479.730 2205.890 1480.910 2207.070 ;
        RECT 1479.730 2204.290 1480.910 2205.470 ;
        RECT 1479.730 2025.890 1480.910 2027.070 ;
        RECT 1479.730 2024.290 1480.910 2025.470 ;
        RECT 1479.730 1845.890 1480.910 1847.070 ;
        RECT 1479.730 1844.290 1480.910 1845.470 ;
        RECT 1479.730 1665.890 1480.910 1667.070 ;
        RECT 1479.730 1664.290 1480.910 1665.470 ;
        RECT 1479.730 1485.890 1480.910 1487.070 ;
        RECT 1479.730 1484.290 1480.910 1485.470 ;
        RECT 1479.730 1305.890 1480.910 1307.070 ;
        RECT 1479.730 1304.290 1480.910 1305.470 ;
        RECT 1479.730 1125.890 1480.910 1127.070 ;
        RECT 1479.730 1124.290 1480.910 1125.470 ;
        RECT 1479.730 945.890 1480.910 947.070 ;
        RECT 1479.730 944.290 1480.910 945.470 ;
        RECT 1479.730 765.890 1480.910 767.070 ;
        RECT 1479.730 764.290 1480.910 765.470 ;
        RECT 1479.730 585.890 1480.910 587.070 ;
        RECT 1479.730 584.290 1480.910 585.470 ;
        RECT 1479.730 405.890 1480.910 407.070 ;
        RECT 1479.730 404.290 1480.910 405.470 ;
        RECT 1479.730 225.890 1480.910 227.070 ;
        RECT 1479.730 224.290 1480.910 225.470 ;
        RECT 1479.730 45.890 1480.910 47.070 ;
        RECT 1479.730 44.290 1480.910 45.470 ;
        RECT 1479.730 -21.310 1480.910 -20.130 ;
        RECT 1479.730 -22.910 1480.910 -21.730 ;
        RECT 1659.730 3541.410 1660.910 3542.590 ;
        RECT 1659.730 3539.810 1660.910 3540.990 ;
        RECT 1659.730 3465.890 1660.910 3467.070 ;
        RECT 1659.730 3464.290 1660.910 3465.470 ;
        RECT 1659.730 3285.890 1660.910 3287.070 ;
        RECT 1659.730 3284.290 1660.910 3285.470 ;
        RECT 1659.730 3105.890 1660.910 3107.070 ;
        RECT 1659.730 3104.290 1660.910 3105.470 ;
        RECT 1659.730 2925.890 1660.910 2927.070 ;
        RECT 1659.730 2924.290 1660.910 2925.470 ;
        RECT 1659.730 2745.890 1660.910 2747.070 ;
        RECT 1659.730 2744.290 1660.910 2745.470 ;
        RECT 1659.730 2565.890 1660.910 2567.070 ;
        RECT 1659.730 2564.290 1660.910 2565.470 ;
        RECT 1659.730 2385.890 1660.910 2387.070 ;
        RECT 1659.730 2384.290 1660.910 2385.470 ;
        RECT 1659.730 2205.890 1660.910 2207.070 ;
        RECT 1659.730 2204.290 1660.910 2205.470 ;
        RECT 1659.730 2025.890 1660.910 2027.070 ;
        RECT 1659.730 2024.290 1660.910 2025.470 ;
        RECT 1659.730 1845.890 1660.910 1847.070 ;
        RECT 1659.730 1844.290 1660.910 1845.470 ;
        RECT 1659.730 1665.890 1660.910 1667.070 ;
        RECT 1659.730 1664.290 1660.910 1665.470 ;
        RECT 1659.730 1485.890 1660.910 1487.070 ;
        RECT 1659.730 1484.290 1660.910 1485.470 ;
        RECT 1659.730 1305.890 1660.910 1307.070 ;
        RECT 1659.730 1304.290 1660.910 1305.470 ;
        RECT 1659.730 1125.890 1660.910 1127.070 ;
        RECT 1659.730 1124.290 1660.910 1125.470 ;
        RECT 1659.730 945.890 1660.910 947.070 ;
        RECT 1659.730 944.290 1660.910 945.470 ;
        RECT 1659.730 765.890 1660.910 767.070 ;
        RECT 1659.730 764.290 1660.910 765.470 ;
        RECT 1659.730 585.890 1660.910 587.070 ;
        RECT 1659.730 584.290 1660.910 585.470 ;
        RECT 1659.730 405.890 1660.910 407.070 ;
        RECT 1659.730 404.290 1660.910 405.470 ;
        RECT 1659.730 225.890 1660.910 227.070 ;
        RECT 1659.730 224.290 1660.910 225.470 ;
        RECT 1659.730 45.890 1660.910 47.070 ;
        RECT 1659.730 44.290 1660.910 45.470 ;
        RECT 1659.730 -21.310 1660.910 -20.130 ;
        RECT 1659.730 -22.910 1660.910 -21.730 ;
        RECT 1839.730 3541.410 1840.910 3542.590 ;
        RECT 1839.730 3539.810 1840.910 3540.990 ;
        RECT 1839.730 3465.890 1840.910 3467.070 ;
        RECT 1839.730 3464.290 1840.910 3465.470 ;
        RECT 1839.730 3285.890 1840.910 3287.070 ;
        RECT 1839.730 3284.290 1840.910 3285.470 ;
        RECT 1839.730 3105.890 1840.910 3107.070 ;
        RECT 1839.730 3104.290 1840.910 3105.470 ;
        RECT 1839.730 2925.890 1840.910 2927.070 ;
        RECT 1839.730 2924.290 1840.910 2925.470 ;
        RECT 1839.730 2745.890 1840.910 2747.070 ;
        RECT 1839.730 2744.290 1840.910 2745.470 ;
        RECT 1839.730 2565.890 1840.910 2567.070 ;
        RECT 1839.730 2564.290 1840.910 2565.470 ;
        RECT 1839.730 2385.890 1840.910 2387.070 ;
        RECT 1839.730 2384.290 1840.910 2385.470 ;
        RECT 1839.730 2205.890 1840.910 2207.070 ;
        RECT 1839.730 2204.290 1840.910 2205.470 ;
        RECT 1839.730 2025.890 1840.910 2027.070 ;
        RECT 1839.730 2024.290 1840.910 2025.470 ;
        RECT 1839.730 1845.890 1840.910 1847.070 ;
        RECT 1839.730 1844.290 1840.910 1845.470 ;
        RECT 1839.730 1665.890 1840.910 1667.070 ;
        RECT 1839.730 1664.290 1840.910 1665.470 ;
        RECT 1839.730 1485.890 1840.910 1487.070 ;
        RECT 1839.730 1484.290 1840.910 1485.470 ;
        RECT 1839.730 1305.890 1840.910 1307.070 ;
        RECT 1839.730 1304.290 1840.910 1305.470 ;
        RECT 1839.730 1125.890 1840.910 1127.070 ;
        RECT 1839.730 1124.290 1840.910 1125.470 ;
        RECT 1839.730 945.890 1840.910 947.070 ;
        RECT 1839.730 944.290 1840.910 945.470 ;
        RECT 1839.730 765.890 1840.910 767.070 ;
        RECT 1839.730 764.290 1840.910 765.470 ;
        RECT 1839.730 585.890 1840.910 587.070 ;
        RECT 1839.730 584.290 1840.910 585.470 ;
        RECT 1839.730 405.890 1840.910 407.070 ;
        RECT 1839.730 404.290 1840.910 405.470 ;
        RECT 1839.730 225.890 1840.910 227.070 ;
        RECT 1839.730 224.290 1840.910 225.470 ;
        RECT 1839.730 45.890 1840.910 47.070 ;
        RECT 1839.730 44.290 1840.910 45.470 ;
        RECT 1839.730 -21.310 1840.910 -20.130 ;
        RECT 1839.730 -22.910 1840.910 -21.730 ;
        RECT 2019.730 3541.410 2020.910 3542.590 ;
        RECT 2019.730 3539.810 2020.910 3540.990 ;
        RECT 2019.730 3465.890 2020.910 3467.070 ;
        RECT 2019.730 3464.290 2020.910 3465.470 ;
        RECT 2019.730 3285.890 2020.910 3287.070 ;
        RECT 2019.730 3284.290 2020.910 3285.470 ;
        RECT 2019.730 3105.890 2020.910 3107.070 ;
        RECT 2019.730 3104.290 2020.910 3105.470 ;
        RECT 2019.730 2925.890 2020.910 2927.070 ;
        RECT 2019.730 2924.290 2020.910 2925.470 ;
        RECT 2019.730 2745.890 2020.910 2747.070 ;
        RECT 2019.730 2744.290 2020.910 2745.470 ;
        RECT 2019.730 2565.890 2020.910 2567.070 ;
        RECT 2019.730 2564.290 2020.910 2565.470 ;
        RECT 2019.730 2385.890 2020.910 2387.070 ;
        RECT 2019.730 2384.290 2020.910 2385.470 ;
        RECT 2019.730 2205.890 2020.910 2207.070 ;
        RECT 2019.730 2204.290 2020.910 2205.470 ;
        RECT 2019.730 2025.890 2020.910 2027.070 ;
        RECT 2019.730 2024.290 2020.910 2025.470 ;
        RECT 2019.730 1845.890 2020.910 1847.070 ;
        RECT 2019.730 1844.290 2020.910 1845.470 ;
        RECT 2019.730 1665.890 2020.910 1667.070 ;
        RECT 2019.730 1664.290 2020.910 1665.470 ;
        RECT 2019.730 1485.890 2020.910 1487.070 ;
        RECT 2019.730 1484.290 2020.910 1485.470 ;
        RECT 2019.730 1305.890 2020.910 1307.070 ;
        RECT 2019.730 1304.290 2020.910 1305.470 ;
        RECT 2019.730 1125.890 2020.910 1127.070 ;
        RECT 2019.730 1124.290 2020.910 1125.470 ;
        RECT 2019.730 945.890 2020.910 947.070 ;
        RECT 2019.730 944.290 2020.910 945.470 ;
        RECT 2019.730 765.890 2020.910 767.070 ;
        RECT 2019.730 764.290 2020.910 765.470 ;
        RECT 2019.730 585.890 2020.910 587.070 ;
        RECT 2019.730 584.290 2020.910 585.470 ;
        RECT 2019.730 405.890 2020.910 407.070 ;
        RECT 2019.730 404.290 2020.910 405.470 ;
        RECT 2019.730 225.890 2020.910 227.070 ;
        RECT 2019.730 224.290 2020.910 225.470 ;
        RECT 2019.730 45.890 2020.910 47.070 ;
        RECT 2019.730 44.290 2020.910 45.470 ;
        RECT 2019.730 -21.310 2020.910 -20.130 ;
        RECT 2019.730 -22.910 2020.910 -21.730 ;
        RECT 2199.730 3541.410 2200.910 3542.590 ;
        RECT 2199.730 3539.810 2200.910 3540.990 ;
        RECT 2199.730 3465.890 2200.910 3467.070 ;
        RECT 2199.730 3464.290 2200.910 3465.470 ;
        RECT 2199.730 3285.890 2200.910 3287.070 ;
        RECT 2199.730 3284.290 2200.910 3285.470 ;
        RECT 2199.730 3105.890 2200.910 3107.070 ;
        RECT 2199.730 3104.290 2200.910 3105.470 ;
        RECT 2199.730 2925.890 2200.910 2927.070 ;
        RECT 2199.730 2924.290 2200.910 2925.470 ;
        RECT 2199.730 2745.890 2200.910 2747.070 ;
        RECT 2199.730 2744.290 2200.910 2745.470 ;
        RECT 2199.730 2565.890 2200.910 2567.070 ;
        RECT 2199.730 2564.290 2200.910 2565.470 ;
        RECT 2199.730 2385.890 2200.910 2387.070 ;
        RECT 2199.730 2384.290 2200.910 2385.470 ;
        RECT 2199.730 2205.890 2200.910 2207.070 ;
        RECT 2199.730 2204.290 2200.910 2205.470 ;
        RECT 2199.730 2025.890 2200.910 2027.070 ;
        RECT 2199.730 2024.290 2200.910 2025.470 ;
        RECT 2199.730 1845.890 2200.910 1847.070 ;
        RECT 2199.730 1844.290 2200.910 1845.470 ;
        RECT 2199.730 1665.890 2200.910 1667.070 ;
        RECT 2199.730 1664.290 2200.910 1665.470 ;
        RECT 2199.730 1485.890 2200.910 1487.070 ;
        RECT 2199.730 1484.290 2200.910 1485.470 ;
        RECT 2199.730 1305.890 2200.910 1307.070 ;
        RECT 2199.730 1304.290 2200.910 1305.470 ;
        RECT 2199.730 1125.890 2200.910 1127.070 ;
        RECT 2199.730 1124.290 2200.910 1125.470 ;
        RECT 2199.730 945.890 2200.910 947.070 ;
        RECT 2199.730 944.290 2200.910 945.470 ;
        RECT 2199.730 765.890 2200.910 767.070 ;
        RECT 2199.730 764.290 2200.910 765.470 ;
        RECT 2199.730 585.890 2200.910 587.070 ;
        RECT 2199.730 584.290 2200.910 585.470 ;
        RECT 2199.730 405.890 2200.910 407.070 ;
        RECT 2199.730 404.290 2200.910 405.470 ;
        RECT 2199.730 225.890 2200.910 227.070 ;
        RECT 2199.730 224.290 2200.910 225.470 ;
        RECT 2199.730 45.890 2200.910 47.070 ;
        RECT 2199.730 44.290 2200.910 45.470 ;
        RECT 2199.730 -21.310 2200.910 -20.130 ;
        RECT 2199.730 -22.910 2200.910 -21.730 ;
        RECT 2379.730 3541.410 2380.910 3542.590 ;
        RECT 2379.730 3539.810 2380.910 3540.990 ;
        RECT 2379.730 3465.890 2380.910 3467.070 ;
        RECT 2379.730 3464.290 2380.910 3465.470 ;
        RECT 2379.730 3285.890 2380.910 3287.070 ;
        RECT 2379.730 3284.290 2380.910 3285.470 ;
        RECT 2379.730 3105.890 2380.910 3107.070 ;
        RECT 2379.730 3104.290 2380.910 3105.470 ;
        RECT 2379.730 2925.890 2380.910 2927.070 ;
        RECT 2379.730 2924.290 2380.910 2925.470 ;
        RECT 2379.730 2745.890 2380.910 2747.070 ;
        RECT 2379.730 2744.290 2380.910 2745.470 ;
        RECT 2379.730 2565.890 2380.910 2567.070 ;
        RECT 2379.730 2564.290 2380.910 2565.470 ;
        RECT 2379.730 2385.890 2380.910 2387.070 ;
        RECT 2379.730 2384.290 2380.910 2385.470 ;
        RECT 2379.730 2205.890 2380.910 2207.070 ;
        RECT 2379.730 2204.290 2380.910 2205.470 ;
        RECT 2379.730 2025.890 2380.910 2027.070 ;
        RECT 2379.730 2024.290 2380.910 2025.470 ;
        RECT 2379.730 1845.890 2380.910 1847.070 ;
        RECT 2379.730 1844.290 2380.910 1845.470 ;
        RECT 2379.730 1665.890 2380.910 1667.070 ;
        RECT 2379.730 1664.290 2380.910 1665.470 ;
        RECT 2379.730 1485.890 2380.910 1487.070 ;
        RECT 2379.730 1484.290 2380.910 1485.470 ;
        RECT 2379.730 1305.890 2380.910 1307.070 ;
        RECT 2379.730 1304.290 2380.910 1305.470 ;
        RECT 2379.730 1125.890 2380.910 1127.070 ;
        RECT 2379.730 1124.290 2380.910 1125.470 ;
        RECT 2379.730 945.890 2380.910 947.070 ;
        RECT 2379.730 944.290 2380.910 945.470 ;
        RECT 2379.730 765.890 2380.910 767.070 ;
        RECT 2379.730 764.290 2380.910 765.470 ;
        RECT 2379.730 585.890 2380.910 587.070 ;
        RECT 2379.730 584.290 2380.910 585.470 ;
        RECT 2379.730 405.890 2380.910 407.070 ;
        RECT 2379.730 404.290 2380.910 405.470 ;
        RECT 2379.730 225.890 2380.910 227.070 ;
        RECT 2379.730 224.290 2380.910 225.470 ;
        RECT 2379.730 45.890 2380.910 47.070 ;
        RECT 2379.730 44.290 2380.910 45.470 ;
        RECT 2379.730 -21.310 2380.910 -20.130 ;
        RECT 2379.730 -22.910 2380.910 -21.730 ;
        RECT 2559.730 3541.410 2560.910 3542.590 ;
        RECT 2559.730 3539.810 2560.910 3540.990 ;
        RECT 2559.730 3465.890 2560.910 3467.070 ;
        RECT 2559.730 3464.290 2560.910 3465.470 ;
        RECT 2559.730 3285.890 2560.910 3287.070 ;
        RECT 2559.730 3284.290 2560.910 3285.470 ;
        RECT 2559.730 3105.890 2560.910 3107.070 ;
        RECT 2559.730 3104.290 2560.910 3105.470 ;
        RECT 2559.730 2925.890 2560.910 2927.070 ;
        RECT 2559.730 2924.290 2560.910 2925.470 ;
        RECT 2559.730 2745.890 2560.910 2747.070 ;
        RECT 2559.730 2744.290 2560.910 2745.470 ;
        RECT 2559.730 2565.890 2560.910 2567.070 ;
        RECT 2559.730 2564.290 2560.910 2565.470 ;
        RECT 2559.730 2385.890 2560.910 2387.070 ;
        RECT 2559.730 2384.290 2560.910 2385.470 ;
        RECT 2559.730 2205.890 2560.910 2207.070 ;
        RECT 2559.730 2204.290 2560.910 2205.470 ;
        RECT 2559.730 2025.890 2560.910 2027.070 ;
        RECT 2559.730 2024.290 2560.910 2025.470 ;
        RECT 2559.730 1845.890 2560.910 1847.070 ;
        RECT 2559.730 1844.290 2560.910 1845.470 ;
        RECT 2559.730 1665.890 2560.910 1667.070 ;
        RECT 2559.730 1664.290 2560.910 1665.470 ;
        RECT 2559.730 1485.890 2560.910 1487.070 ;
        RECT 2559.730 1484.290 2560.910 1485.470 ;
        RECT 2559.730 1305.890 2560.910 1307.070 ;
        RECT 2559.730 1304.290 2560.910 1305.470 ;
        RECT 2559.730 1125.890 2560.910 1127.070 ;
        RECT 2559.730 1124.290 2560.910 1125.470 ;
        RECT 2559.730 945.890 2560.910 947.070 ;
        RECT 2559.730 944.290 2560.910 945.470 ;
        RECT 2559.730 765.890 2560.910 767.070 ;
        RECT 2559.730 764.290 2560.910 765.470 ;
        RECT 2559.730 585.890 2560.910 587.070 ;
        RECT 2559.730 584.290 2560.910 585.470 ;
        RECT 2559.730 405.890 2560.910 407.070 ;
        RECT 2559.730 404.290 2560.910 405.470 ;
        RECT 2559.730 225.890 2560.910 227.070 ;
        RECT 2559.730 224.290 2560.910 225.470 ;
        RECT 2559.730 45.890 2560.910 47.070 ;
        RECT 2559.730 44.290 2560.910 45.470 ;
        RECT 2559.730 -21.310 2560.910 -20.130 ;
        RECT 2559.730 -22.910 2560.910 -21.730 ;
        RECT 2739.730 3541.410 2740.910 3542.590 ;
        RECT 2739.730 3539.810 2740.910 3540.990 ;
        RECT 2739.730 3465.890 2740.910 3467.070 ;
        RECT 2739.730 3464.290 2740.910 3465.470 ;
        RECT 2739.730 3285.890 2740.910 3287.070 ;
        RECT 2739.730 3284.290 2740.910 3285.470 ;
        RECT 2739.730 3105.890 2740.910 3107.070 ;
        RECT 2739.730 3104.290 2740.910 3105.470 ;
        RECT 2739.730 2925.890 2740.910 2927.070 ;
        RECT 2739.730 2924.290 2740.910 2925.470 ;
        RECT 2739.730 2745.890 2740.910 2747.070 ;
        RECT 2739.730 2744.290 2740.910 2745.470 ;
        RECT 2739.730 2565.890 2740.910 2567.070 ;
        RECT 2739.730 2564.290 2740.910 2565.470 ;
        RECT 2739.730 2385.890 2740.910 2387.070 ;
        RECT 2739.730 2384.290 2740.910 2385.470 ;
        RECT 2739.730 2205.890 2740.910 2207.070 ;
        RECT 2739.730 2204.290 2740.910 2205.470 ;
        RECT 2739.730 2025.890 2740.910 2027.070 ;
        RECT 2739.730 2024.290 2740.910 2025.470 ;
        RECT 2739.730 1845.890 2740.910 1847.070 ;
        RECT 2739.730 1844.290 2740.910 1845.470 ;
        RECT 2739.730 1665.890 2740.910 1667.070 ;
        RECT 2739.730 1664.290 2740.910 1665.470 ;
        RECT 2739.730 1485.890 2740.910 1487.070 ;
        RECT 2739.730 1484.290 2740.910 1485.470 ;
        RECT 2739.730 1305.890 2740.910 1307.070 ;
        RECT 2739.730 1304.290 2740.910 1305.470 ;
        RECT 2739.730 1125.890 2740.910 1127.070 ;
        RECT 2739.730 1124.290 2740.910 1125.470 ;
        RECT 2739.730 945.890 2740.910 947.070 ;
        RECT 2739.730 944.290 2740.910 945.470 ;
        RECT 2739.730 765.890 2740.910 767.070 ;
        RECT 2739.730 764.290 2740.910 765.470 ;
        RECT 2739.730 585.890 2740.910 587.070 ;
        RECT 2739.730 584.290 2740.910 585.470 ;
        RECT 2739.730 405.890 2740.910 407.070 ;
        RECT 2739.730 404.290 2740.910 405.470 ;
        RECT 2739.730 225.890 2740.910 227.070 ;
        RECT 2739.730 224.290 2740.910 225.470 ;
        RECT 2739.730 45.890 2740.910 47.070 ;
        RECT 2739.730 44.290 2740.910 45.470 ;
        RECT 2739.730 -21.310 2740.910 -20.130 ;
        RECT 2739.730 -22.910 2740.910 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3465.890 2947.090 3467.070 ;
        RECT 2945.910 3464.290 2947.090 3465.470 ;
        RECT 2945.910 3285.890 2947.090 3287.070 ;
        RECT 2945.910 3284.290 2947.090 3285.470 ;
        RECT 2945.910 3105.890 2947.090 3107.070 ;
        RECT 2945.910 3104.290 2947.090 3105.470 ;
        RECT 2945.910 2925.890 2947.090 2927.070 ;
        RECT 2945.910 2924.290 2947.090 2925.470 ;
        RECT 2945.910 2745.890 2947.090 2747.070 ;
        RECT 2945.910 2744.290 2947.090 2745.470 ;
        RECT 2945.910 2565.890 2947.090 2567.070 ;
        RECT 2945.910 2564.290 2947.090 2565.470 ;
        RECT 2945.910 2385.890 2947.090 2387.070 ;
        RECT 2945.910 2384.290 2947.090 2385.470 ;
        RECT 2945.910 2205.890 2947.090 2207.070 ;
        RECT 2945.910 2204.290 2947.090 2205.470 ;
        RECT 2945.910 2025.890 2947.090 2027.070 ;
        RECT 2945.910 2024.290 2947.090 2025.470 ;
        RECT 2945.910 1845.890 2947.090 1847.070 ;
        RECT 2945.910 1844.290 2947.090 1845.470 ;
        RECT 2945.910 1665.890 2947.090 1667.070 ;
        RECT 2945.910 1664.290 2947.090 1665.470 ;
        RECT 2945.910 1485.890 2947.090 1487.070 ;
        RECT 2945.910 1484.290 2947.090 1485.470 ;
        RECT 2945.910 1305.890 2947.090 1307.070 ;
        RECT 2945.910 1304.290 2947.090 1305.470 ;
        RECT 2945.910 1125.890 2947.090 1127.070 ;
        RECT 2945.910 1124.290 2947.090 1125.470 ;
        RECT 2945.910 945.890 2947.090 947.070 ;
        RECT 2945.910 944.290 2947.090 945.470 ;
        RECT 2945.910 765.890 2947.090 767.070 ;
        RECT 2945.910 764.290 2947.090 765.470 ;
        RECT 2945.910 585.890 2947.090 587.070 ;
        RECT 2945.910 584.290 2947.090 585.470 ;
        RECT 2945.910 405.890 2947.090 407.070 ;
        RECT 2945.910 404.290 2947.090 405.470 ;
        RECT 2945.910 225.890 2947.090 227.070 ;
        RECT 2945.910 224.290 2947.090 225.470 ;
        RECT 2945.910 45.890 2947.090 47.070 ;
        RECT 2945.910 44.290 2947.090 45.470 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.330 3542.650 -25.430 3542.710 ;
        RECT 38.870 3542.650 41.770 3542.710 ;
        RECT 218.870 3542.650 221.770 3542.710 ;
        RECT 398.870 3542.650 401.770 3542.710 ;
        RECT 578.870 3542.650 581.770 3542.710 ;
        RECT 758.870 3542.650 761.770 3542.710 ;
        RECT 938.870 3542.650 941.770 3542.710 ;
        RECT 1118.870 3542.650 1121.770 3542.710 ;
        RECT 1298.870 3542.650 1301.770 3542.710 ;
        RECT 1478.870 3542.650 1481.770 3542.710 ;
        RECT 1658.870 3542.650 1661.770 3542.710 ;
        RECT 1838.870 3542.650 1841.770 3542.710 ;
        RECT 2018.870 3542.650 2021.770 3542.710 ;
        RECT 2198.870 3542.650 2201.770 3542.710 ;
        RECT 2378.870 3542.650 2381.770 3542.710 ;
        RECT 2558.870 3542.650 2561.770 3542.710 ;
        RECT 2738.870 3542.650 2741.770 3542.710 ;
        RECT 2945.050 3542.650 2947.950 3542.710 ;
        RECT -28.330 3539.750 2947.950 3542.650 ;
        RECT -28.330 3539.690 -25.430 3539.750 ;
        RECT 38.870 3539.690 41.770 3539.750 ;
        RECT 218.870 3539.690 221.770 3539.750 ;
        RECT 398.870 3539.690 401.770 3539.750 ;
        RECT 578.870 3539.690 581.770 3539.750 ;
        RECT 758.870 3539.690 761.770 3539.750 ;
        RECT 938.870 3539.690 941.770 3539.750 ;
        RECT 1118.870 3539.690 1121.770 3539.750 ;
        RECT 1298.870 3539.690 1301.770 3539.750 ;
        RECT 1478.870 3539.690 1481.770 3539.750 ;
        RECT 1658.870 3539.690 1661.770 3539.750 ;
        RECT 1838.870 3539.690 1841.770 3539.750 ;
        RECT 2018.870 3539.690 2021.770 3539.750 ;
        RECT 2198.870 3539.690 2201.770 3539.750 ;
        RECT 2378.870 3539.690 2381.770 3539.750 ;
        RECT 2558.870 3539.690 2561.770 3539.750 ;
        RECT 2738.870 3539.690 2741.770 3539.750 ;
        RECT 2945.050 3539.690 2947.950 3539.750 ;
        RECT -28.330 3467.130 -25.430 3467.190 ;
        RECT 38.870 3467.130 41.770 3467.190 ;
        RECT 218.870 3467.130 221.770 3467.190 ;
        RECT 398.870 3467.130 401.770 3467.190 ;
        RECT 578.870 3467.130 581.770 3467.190 ;
        RECT 758.870 3467.130 761.770 3467.190 ;
        RECT 938.870 3467.130 941.770 3467.190 ;
        RECT 1118.870 3467.130 1121.770 3467.190 ;
        RECT 1298.870 3467.130 1301.770 3467.190 ;
        RECT 1478.870 3467.130 1481.770 3467.190 ;
        RECT 1658.870 3467.130 1661.770 3467.190 ;
        RECT 1838.870 3467.130 1841.770 3467.190 ;
        RECT 2018.870 3467.130 2021.770 3467.190 ;
        RECT 2198.870 3467.130 2201.770 3467.190 ;
        RECT 2378.870 3467.130 2381.770 3467.190 ;
        RECT 2558.870 3467.130 2561.770 3467.190 ;
        RECT 2738.870 3467.130 2741.770 3467.190 ;
        RECT 2945.050 3467.130 2947.950 3467.190 ;
        RECT -32.930 3464.230 2952.550 3467.130 ;
        RECT -28.330 3464.170 -25.430 3464.230 ;
        RECT 38.870 3464.170 41.770 3464.230 ;
        RECT 218.870 3464.170 221.770 3464.230 ;
        RECT 398.870 3464.170 401.770 3464.230 ;
        RECT 578.870 3464.170 581.770 3464.230 ;
        RECT 758.870 3464.170 761.770 3464.230 ;
        RECT 938.870 3464.170 941.770 3464.230 ;
        RECT 1118.870 3464.170 1121.770 3464.230 ;
        RECT 1298.870 3464.170 1301.770 3464.230 ;
        RECT 1478.870 3464.170 1481.770 3464.230 ;
        RECT 1658.870 3464.170 1661.770 3464.230 ;
        RECT 1838.870 3464.170 1841.770 3464.230 ;
        RECT 2018.870 3464.170 2021.770 3464.230 ;
        RECT 2198.870 3464.170 2201.770 3464.230 ;
        RECT 2378.870 3464.170 2381.770 3464.230 ;
        RECT 2558.870 3464.170 2561.770 3464.230 ;
        RECT 2738.870 3464.170 2741.770 3464.230 ;
        RECT 2945.050 3464.170 2947.950 3464.230 ;
        RECT -28.330 3287.130 -25.430 3287.190 ;
        RECT 38.870 3287.130 41.770 3287.190 ;
        RECT 218.870 3287.130 221.770 3287.190 ;
        RECT 398.870 3287.130 401.770 3287.190 ;
        RECT 578.870 3287.130 581.770 3287.190 ;
        RECT 758.870 3287.130 761.770 3287.190 ;
        RECT 938.870 3287.130 941.770 3287.190 ;
        RECT 1118.870 3287.130 1121.770 3287.190 ;
        RECT 1298.870 3287.130 1301.770 3287.190 ;
        RECT 1478.870 3287.130 1481.770 3287.190 ;
        RECT 1658.870 3287.130 1661.770 3287.190 ;
        RECT 1838.870 3287.130 1841.770 3287.190 ;
        RECT 2018.870 3287.130 2021.770 3287.190 ;
        RECT 2198.870 3287.130 2201.770 3287.190 ;
        RECT 2378.870 3287.130 2381.770 3287.190 ;
        RECT 2558.870 3287.130 2561.770 3287.190 ;
        RECT 2738.870 3287.130 2741.770 3287.190 ;
        RECT 2945.050 3287.130 2947.950 3287.190 ;
        RECT -32.930 3284.230 2952.550 3287.130 ;
        RECT -28.330 3284.170 -25.430 3284.230 ;
        RECT 38.870 3284.170 41.770 3284.230 ;
        RECT 218.870 3284.170 221.770 3284.230 ;
        RECT 398.870 3284.170 401.770 3284.230 ;
        RECT 578.870 3284.170 581.770 3284.230 ;
        RECT 758.870 3284.170 761.770 3284.230 ;
        RECT 938.870 3284.170 941.770 3284.230 ;
        RECT 1118.870 3284.170 1121.770 3284.230 ;
        RECT 1298.870 3284.170 1301.770 3284.230 ;
        RECT 1478.870 3284.170 1481.770 3284.230 ;
        RECT 1658.870 3284.170 1661.770 3284.230 ;
        RECT 1838.870 3284.170 1841.770 3284.230 ;
        RECT 2018.870 3284.170 2021.770 3284.230 ;
        RECT 2198.870 3284.170 2201.770 3284.230 ;
        RECT 2378.870 3284.170 2381.770 3284.230 ;
        RECT 2558.870 3284.170 2561.770 3284.230 ;
        RECT 2738.870 3284.170 2741.770 3284.230 ;
        RECT 2945.050 3284.170 2947.950 3284.230 ;
        RECT -28.330 3107.130 -25.430 3107.190 ;
        RECT 38.870 3107.130 41.770 3107.190 ;
        RECT 218.870 3107.130 221.770 3107.190 ;
        RECT 398.870 3107.130 401.770 3107.190 ;
        RECT 578.870 3107.130 581.770 3107.190 ;
        RECT 758.870 3107.130 761.770 3107.190 ;
        RECT 938.870 3107.130 941.770 3107.190 ;
        RECT 1118.870 3107.130 1121.770 3107.190 ;
        RECT 1298.870 3107.130 1301.770 3107.190 ;
        RECT 1478.870 3107.130 1481.770 3107.190 ;
        RECT 1658.870 3107.130 1661.770 3107.190 ;
        RECT 1838.870 3107.130 1841.770 3107.190 ;
        RECT 2018.870 3107.130 2021.770 3107.190 ;
        RECT 2198.870 3107.130 2201.770 3107.190 ;
        RECT 2378.870 3107.130 2381.770 3107.190 ;
        RECT 2558.870 3107.130 2561.770 3107.190 ;
        RECT 2738.870 3107.130 2741.770 3107.190 ;
        RECT 2945.050 3107.130 2947.950 3107.190 ;
        RECT -32.930 3104.230 2952.550 3107.130 ;
        RECT -28.330 3104.170 -25.430 3104.230 ;
        RECT 38.870 3104.170 41.770 3104.230 ;
        RECT 218.870 3104.170 221.770 3104.230 ;
        RECT 398.870 3104.170 401.770 3104.230 ;
        RECT 578.870 3104.170 581.770 3104.230 ;
        RECT 758.870 3104.170 761.770 3104.230 ;
        RECT 938.870 3104.170 941.770 3104.230 ;
        RECT 1118.870 3104.170 1121.770 3104.230 ;
        RECT 1298.870 3104.170 1301.770 3104.230 ;
        RECT 1478.870 3104.170 1481.770 3104.230 ;
        RECT 1658.870 3104.170 1661.770 3104.230 ;
        RECT 1838.870 3104.170 1841.770 3104.230 ;
        RECT 2018.870 3104.170 2021.770 3104.230 ;
        RECT 2198.870 3104.170 2201.770 3104.230 ;
        RECT 2378.870 3104.170 2381.770 3104.230 ;
        RECT 2558.870 3104.170 2561.770 3104.230 ;
        RECT 2738.870 3104.170 2741.770 3104.230 ;
        RECT 2945.050 3104.170 2947.950 3104.230 ;
        RECT -28.330 2927.130 -25.430 2927.190 ;
        RECT 38.870 2927.130 41.770 2927.190 ;
        RECT 218.870 2927.130 221.770 2927.190 ;
        RECT 398.870 2927.130 401.770 2927.190 ;
        RECT 578.870 2927.130 581.770 2927.190 ;
        RECT 758.870 2927.130 761.770 2927.190 ;
        RECT 938.870 2927.130 941.770 2927.190 ;
        RECT 1118.870 2927.130 1121.770 2927.190 ;
        RECT 1298.870 2927.130 1301.770 2927.190 ;
        RECT 1478.870 2927.130 1481.770 2927.190 ;
        RECT 1658.870 2927.130 1661.770 2927.190 ;
        RECT 1838.870 2927.130 1841.770 2927.190 ;
        RECT 2018.870 2927.130 2021.770 2927.190 ;
        RECT 2198.870 2927.130 2201.770 2927.190 ;
        RECT 2378.870 2927.130 2381.770 2927.190 ;
        RECT 2558.870 2927.130 2561.770 2927.190 ;
        RECT 2738.870 2927.130 2741.770 2927.190 ;
        RECT 2945.050 2927.130 2947.950 2927.190 ;
        RECT -32.930 2924.230 2952.550 2927.130 ;
        RECT -28.330 2924.170 -25.430 2924.230 ;
        RECT 38.870 2924.170 41.770 2924.230 ;
        RECT 218.870 2924.170 221.770 2924.230 ;
        RECT 398.870 2924.170 401.770 2924.230 ;
        RECT 578.870 2924.170 581.770 2924.230 ;
        RECT 758.870 2924.170 761.770 2924.230 ;
        RECT 938.870 2924.170 941.770 2924.230 ;
        RECT 1118.870 2924.170 1121.770 2924.230 ;
        RECT 1298.870 2924.170 1301.770 2924.230 ;
        RECT 1478.870 2924.170 1481.770 2924.230 ;
        RECT 1658.870 2924.170 1661.770 2924.230 ;
        RECT 1838.870 2924.170 1841.770 2924.230 ;
        RECT 2018.870 2924.170 2021.770 2924.230 ;
        RECT 2198.870 2924.170 2201.770 2924.230 ;
        RECT 2378.870 2924.170 2381.770 2924.230 ;
        RECT 2558.870 2924.170 2561.770 2924.230 ;
        RECT 2738.870 2924.170 2741.770 2924.230 ;
        RECT 2945.050 2924.170 2947.950 2924.230 ;
        RECT -28.330 2747.130 -25.430 2747.190 ;
        RECT 38.870 2747.130 41.770 2747.190 ;
        RECT 218.870 2747.130 221.770 2747.190 ;
        RECT 398.870 2747.130 401.770 2747.190 ;
        RECT 578.870 2747.130 581.770 2747.190 ;
        RECT 758.870 2747.130 761.770 2747.190 ;
        RECT 938.870 2747.130 941.770 2747.190 ;
        RECT 1118.870 2747.130 1121.770 2747.190 ;
        RECT 1298.870 2747.130 1301.770 2747.190 ;
        RECT 1478.870 2747.130 1481.770 2747.190 ;
        RECT 1658.870 2747.130 1661.770 2747.190 ;
        RECT 1838.870 2747.130 1841.770 2747.190 ;
        RECT 2018.870 2747.130 2021.770 2747.190 ;
        RECT 2198.870 2747.130 2201.770 2747.190 ;
        RECT 2378.870 2747.130 2381.770 2747.190 ;
        RECT 2558.870 2747.130 2561.770 2747.190 ;
        RECT 2738.870 2747.130 2741.770 2747.190 ;
        RECT 2945.050 2747.130 2947.950 2747.190 ;
        RECT -32.930 2744.230 2952.550 2747.130 ;
        RECT -28.330 2744.170 -25.430 2744.230 ;
        RECT 38.870 2744.170 41.770 2744.230 ;
        RECT 218.870 2744.170 221.770 2744.230 ;
        RECT 398.870 2744.170 401.770 2744.230 ;
        RECT 578.870 2744.170 581.770 2744.230 ;
        RECT 758.870 2744.170 761.770 2744.230 ;
        RECT 938.870 2744.170 941.770 2744.230 ;
        RECT 1118.870 2744.170 1121.770 2744.230 ;
        RECT 1298.870 2744.170 1301.770 2744.230 ;
        RECT 1478.870 2744.170 1481.770 2744.230 ;
        RECT 1658.870 2744.170 1661.770 2744.230 ;
        RECT 1838.870 2744.170 1841.770 2744.230 ;
        RECT 2018.870 2744.170 2021.770 2744.230 ;
        RECT 2198.870 2744.170 2201.770 2744.230 ;
        RECT 2378.870 2744.170 2381.770 2744.230 ;
        RECT 2558.870 2744.170 2561.770 2744.230 ;
        RECT 2738.870 2744.170 2741.770 2744.230 ;
        RECT 2945.050 2744.170 2947.950 2744.230 ;
        RECT -28.330 2567.130 -25.430 2567.190 ;
        RECT 38.870 2567.130 41.770 2567.190 ;
        RECT 218.870 2567.130 221.770 2567.190 ;
        RECT 398.870 2567.130 401.770 2567.190 ;
        RECT 578.870 2567.130 581.770 2567.190 ;
        RECT 758.870 2567.130 761.770 2567.190 ;
        RECT 938.870 2567.130 941.770 2567.190 ;
        RECT 1118.870 2567.130 1121.770 2567.190 ;
        RECT 1298.870 2567.130 1301.770 2567.190 ;
        RECT 1478.870 2567.130 1481.770 2567.190 ;
        RECT 1658.870 2567.130 1661.770 2567.190 ;
        RECT 1838.870 2567.130 1841.770 2567.190 ;
        RECT 2018.870 2567.130 2021.770 2567.190 ;
        RECT 2198.870 2567.130 2201.770 2567.190 ;
        RECT 2378.870 2567.130 2381.770 2567.190 ;
        RECT 2558.870 2567.130 2561.770 2567.190 ;
        RECT 2738.870 2567.130 2741.770 2567.190 ;
        RECT 2945.050 2567.130 2947.950 2567.190 ;
        RECT -32.930 2564.230 2952.550 2567.130 ;
        RECT -28.330 2564.170 -25.430 2564.230 ;
        RECT 38.870 2564.170 41.770 2564.230 ;
        RECT 218.870 2564.170 221.770 2564.230 ;
        RECT 398.870 2564.170 401.770 2564.230 ;
        RECT 578.870 2564.170 581.770 2564.230 ;
        RECT 758.870 2564.170 761.770 2564.230 ;
        RECT 938.870 2564.170 941.770 2564.230 ;
        RECT 1118.870 2564.170 1121.770 2564.230 ;
        RECT 1298.870 2564.170 1301.770 2564.230 ;
        RECT 1478.870 2564.170 1481.770 2564.230 ;
        RECT 1658.870 2564.170 1661.770 2564.230 ;
        RECT 1838.870 2564.170 1841.770 2564.230 ;
        RECT 2018.870 2564.170 2021.770 2564.230 ;
        RECT 2198.870 2564.170 2201.770 2564.230 ;
        RECT 2378.870 2564.170 2381.770 2564.230 ;
        RECT 2558.870 2564.170 2561.770 2564.230 ;
        RECT 2738.870 2564.170 2741.770 2564.230 ;
        RECT 2945.050 2564.170 2947.950 2564.230 ;
        RECT -28.330 2387.130 -25.430 2387.190 ;
        RECT 38.870 2387.130 41.770 2387.190 ;
        RECT 218.870 2387.130 221.770 2387.190 ;
        RECT 398.870 2387.130 401.770 2387.190 ;
        RECT 578.870 2387.130 581.770 2387.190 ;
        RECT 758.870 2387.130 761.770 2387.190 ;
        RECT 938.870 2387.130 941.770 2387.190 ;
        RECT 1118.870 2387.130 1121.770 2387.190 ;
        RECT 1298.870 2387.130 1301.770 2387.190 ;
        RECT 1478.870 2387.130 1481.770 2387.190 ;
        RECT 1658.870 2387.130 1661.770 2387.190 ;
        RECT 1838.870 2387.130 1841.770 2387.190 ;
        RECT 2018.870 2387.130 2021.770 2387.190 ;
        RECT 2198.870 2387.130 2201.770 2387.190 ;
        RECT 2378.870 2387.130 2381.770 2387.190 ;
        RECT 2558.870 2387.130 2561.770 2387.190 ;
        RECT 2738.870 2387.130 2741.770 2387.190 ;
        RECT 2945.050 2387.130 2947.950 2387.190 ;
        RECT -32.930 2384.230 2952.550 2387.130 ;
        RECT -28.330 2384.170 -25.430 2384.230 ;
        RECT 38.870 2384.170 41.770 2384.230 ;
        RECT 218.870 2384.170 221.770 2384.230 ;
        RECT 398.870 2384.170 401.770 2384.230 ;
        RECT 578.870 2384.170 581.770 2384.230 ;
        RECT 758.870 2384.170 761.770 2384.230 ;
        RECT 938.870 2384.170 941.770 2384.230 ;
        RECT 1118.870 2384.170 1121.770 2384.230 ;
        RECT 1298.870 2384.170 1301.770 2384.230 ;
        RECT 1478.870 2384.170 1481.770 2384.230 ;
        RECT 1658.870 2384.170 1661.770 2384.230 ;
        RECT 1838.870 2384.170 1841.770 2384.230 ;
        RECT 2018.870 2384.170 2021.770 2384.230 ;
        RECT 2198.870 2384.170 2201.770 2384.230 ;
        RECT 2378.870 2384.170 2381.770 2384.230 ;
        RECT 2558.870 2384.170 2561.770 2384.230 ;
        RECT 2738.870 2384.170 2741.770 2384.230 ;
        RECT 2945.050 2384.170 2947.950 2384.230 ;
        RECT -28.330 2207.130 -25.430 2207.190 ;
        RECT 38.870 2207.130 41.770 2207.190 ;
        RECT 218.870 2207.130 221.770 2207.190 ;
        RECT 398.870 2207.130 401.770 2207.190 ;
        RECT 578.870 2207.130 581.770 2207.190 ;
        RECT 758.870 2207.130 761.770 2207.190 ;
        RECT 938.870 2207.130 941.770 2207.190 ;
        RECT 1118.870 2207.130 1121.770 2207.190 ;
        RECT 1298.870 2207.130 1301.770 2207.190 ;
        RECT 1478.870 2207.130 1481.770 2207.190 ;
        RECT 1658.870 2207.130 1661.770 2207.190 ;
        RECT 1838.870 2207.130 1841.770 2207.190 ;
        RECT 2018.870 2207.130 2021.770 2207.190 ;
        RECT 2198.870 2207.130 2201.770 2207.190 ;
        RECT 2378.870 2207.130 2381.770 2207.190 ;
        RECT 2558.870 2207.130 2561.770 2207.190 ;
        RECT 2738.870 2207.130 2741.770 2207.190 ;
        RECT 2945.050 2207.130 2947.950 2207.190 ;
        RECT -32.930 2204.230 2952.550 2207.130 ;
        RECT -28.330 2204.170 -25.430 2204.230 ;
        RECT 38.870 2204.170 41.770 2204.230 ;
        RECT 218.870 2204.170 221.770 2204.230 ;
        RECT 398.870 2204.170 401.770 2204.230 ;
        RECT 578.870 2204.170 581.770 2204.230 ;
        RECT 758.870 2204.170 761.770 2204.230 ;
        RECT 938.870 2204.170 941.770 2204.230 ;
        RECT 1118.870 2204.170 1121.770 2204.230 ;
        RECT 1298.870 2204.170 1301.770 2204.230 ;
        RECT 1478.870 2204.170 1481.770 2204.230 ;
        RECT 1658.870 2204.170 1661.770 2204.230 ;
        RECT 1838.870 2204.170 1841.770 2204.230 ;
        RECT 2018.870 2204.170 2021.770 2204.230 ;
        RECT 2198.870 2204.170 2201.770 2204.230 ;
        RECT 2378.870 2204.170 2381.770 2204.230 ;
        RECT 2558.870 2204.170 2561.770 2204.230 ;
        RECT 2738.870 2204.170 2741.770 2204.230 ;
        RECT 2945.050 2204.170 2947.950 2204.230 ;
        RECT -28.330 2027.130 -25.430 2027.190 ;
        RECT 38.870 2027.130 41.770 2027.190 ;
        RECT 218.870 2027.130 221.770 2027.190 ;
        RECT 398.870 2027.130 401.770 2027.190 ;
        RECT 578.870 2027.130 581.770 2027.190 ;
        RECT 758.870 2027.130 761.770 2027.190 ;
        RECT 938.870 2027.130 941.770 2027.190 ;
        RECT 1118.870 2027.130 1121.770 2027.190 ;
        RECT 1298.870 2027.130 1301.770 2027.190 ;
        RECT 1478.870 2027.130 1481.770 2027.190 ;
        RECT 1658.870 2027.130 1661.770 2027.190 ;
        RECT 1838.870 2027.130 1841.770 2027.190 ;
        RECT 2018.870 2027.130 2021.770 2027.190 ;
        RECT 2198.870 2027.130 2201.770 2027.190 ;
        RECT 2378.870 2027.130 2381.770 2027.190 ;
        RECT 2558.870 2027.130 2561.770 2027.190 ;
        RECT 2738.870 2027.130 2741.770 2027.190 ;
        RECT 2945.050 2027.130 2947.950 2027.190 ;
        RECT -32.930 2024.230 2952.550 2027.130 ;
        RECT -28.330 2024.170 -25.430 2024.230 ;
        RECT 38.870 2024.170 41.770 2024.230 ;
        RECT 218.870 2024.170 221.770 2024.230 ;
        RECT 398.870 2024.170 401.770 2024.230 ;
        RECT 578.870 2024.170 581.770 2024.230 ;
        RECT 758.870 2024.170 761.770 2024.230 ;
        RECT 938.870 2024.170 941.770 2024.230 ;
        RECT 1118.870 2024.170 1121.770 2024.230 ;
        RECT 1298.870 2024.170 1301.770 2024.230 ;
        RECT 1478.870 2024.170 1481.770 2024.230 ;
        RECT 1658.870 2024.170 1661.770 2024.230 ;
        RECT 1838.870 2024.170 1841.770 2024.230 ;
        RECT 2018.870 2024.170 2021.770 2024.230 ;
        RECT 2198.870 2024.170 2201.770 2024.230 ;
        RECT 2378.870 2024.170 2381.770 2024.230 ;
        RECT 2558.870 2024.170 2561.770 2024.230 ;
        RECT 2738.870 2024.170 2741.770 2024.230 ;
        RECT 2945.050 2024.170 2947.950 2024.230 ;
        RECT -28.330 1847.130 -25.430 1847.190 ;
        RECT 38.870 1847.130 41.770 1847.190 ;
        RECT 218.870 1847.130 221.770 1847.190 ;
        RECT 398.870 1847.130 401.770 1847.190 ;
        RECT 578.870 1847.130 581.770 1847.190 ;
        RECT 758.870 1847.130 761.770 1847.190 ;
        RECT 938.870 1847.130 941.770 1847.190 ;
        RECT 1118.870 1847.130 1121.770 1847.190 ;
        RECT 1298.870 1847.130 1301.770 1847.190 ;
        RECT 1478.870 1847.130 1481.770 1847.190 ;
        RECT 1658.870 1847.130 1661.770 1847.190 ;
        RECT 1838.870 1847.130 1841.770 1847.190 ;
        RECT 2018.870 1847.130 2021.770 1847.190 ;
        RECT 2198.870 1847.130 2201.770 1847.190 ;
        RECT 2378.870 1847.130 2381.770 1847.190 ;
        RECT 2558.870 1847.130 2561.770 1847.190 ;
        RECT 2738.870 1847.130 2741.770 1847.190 ;
        RECT 2945.050 1847.130 2947.950 1847.190 ;
        RECT -32.930 1844.230 2952.550 1847.130 ;
        RECT -28.330 1844.170 -25.430 1844.230 ;
        RECT 38.870 1844.170 41.770 1844.230 ;
        RECT 218.870 1844.170 221.770 1844.230 ;
        RECT 398.870 1844.170 401.770 1844.230 ;
        RECT 578.870 1844.170 581.770 1844.230 ;
        RECT 758.870 1844.170 761.770 1844.230 ;
        RECT 938.870 1844.170 941.770 1844.230 ;
        RECT 1118.870 1844.170 1121.770 1844.230 ;
        RECT 1298.870 1844.170 1301.770 1844.230 ;
        RECT 1478.870 1844.170 1481.770 1844.230 ;
        RECT 1658.870 1844.170 1661.770 1844.230 ;
        RECT 1838.870 1844.170 1841.770 1844.230 ;
        RECT 2018.870 1844.170 2021.770 1844.230 ;
        RECT 2198.870 1844.170 2201.770 1844.230 ;
        RECT 2378.870 1844.170 2381.770 1844.230 ;
        RECT 2558.870 1844.170 2561.770 1844.230 ;
        RECT 2738.870 1844.170 2741.770 1844.230 ;
        RECT 2945.050 1844.170 2947.950 1844.230 ;
        RECT -28.330 1667.130 -25.430 1667.190 ;
        RECT 38.870 1667.130 41.770 1667.190 ;
        RECT 218.870 1667.130 221.770 1667.190 ;
        RECT 398.870 1667.130 401.770 1667.190 ;
        RECT 578.870 1667.130 581.770 1667.190 ;
        RECT 758.870 1667.130 761.770 1667.190 ;
        RECT 938.870 1667.130 941.770 1667.190 ;
        RECT 1118.870 1667.130 1121.770 1667.190 ;
        RECT 1298.870 1667.130 1301.770 1667.190 ;
        RECT 1478.870 1667.130 1481.770 1667.190 ;
        RECT 1658.870 1667.130 1661.770 1667.190 ;
        RECT 1838.870 1667.130 1841.770 1667.190 ;
        RECT 2018.870 1667.130 2021.770 1667.190 ;
        RECT 2198.870 1667.130 2201.770 1667.190 ;
        RECT 2378.870 1667.130 2381.770 1667.190 ;
        RECT 2558.870 1667.130 2561.770 1667.190 ;
        RECT 2738.870 1667.130 2741.770 1667.190 ;
        RECT 2945.050 1667.130 2947.950 1667.190 ;
        RECT -32.930 1664.230 2952.550 1667.130 ;
        RECT -28.330 1664.170 -25.430 1664.230 ;
        RECT 38.870 1664.170 41.770 1664.230 ;
        RECT 218.870 1664.170 221.770 1664.230 ;
        RECT 398.870 1664.170 401.770 1664.230 ;
        RECT 578.870 1664.170 581.770 1664.230 ;
        RECT 758.870 1664.170 761.770 1664.230 ;
        RECT 938.870 1664.170 941.770 1664.230 ;
        RECT 1118.870 1664.170 1121.770 1664.230 ;
        RECT 1298.870 1664.170 1301.770 1664.230 ;
        RECT 1478.870 1664.170 1481.770 1664.230 ;
        RECT 1658.870 1664.170 1661.770 1664.230 ;
        RECT 1838.870 1664.170 1841.770 1664.230 ;
        RECT 2018.870 1664.170 2021.770 1664.230 ;
        RECT 2198.870 1664.170 2201.770 1664.230 ;
        RECT 2378.870 1664.170 2381.770 1664.230 ;
        RECT 2558.870 1664.170 2561.770 1664.230 ;
        RECT 2738.870 1664.170 2741.770 1664.230 ;
        RECT 2945.050 1664.170 2947.950 1664.230 ;
        RECT -28.330 1487.130 -25.430 1487.190 ;
        RECT 38.870 1487.130 41.770 1487.190 ;
        RECT 218.870 1487.130 221.770 1487.190 ;
        RECT 398.870 1487.130 401.770 1487.190 ;
        RECT 578.870 1487.130 581.770 1487.190 ;
        RECT 758.870 1487.130 761.770 1487.190 ;
        RECT 938.870 1487.130 941.770 1487.190 ;
        RECT 1118.870 1487.130 1121.770 1487.190 ;
        RECT 1298.870 1487.130 1301.770 1487.190 ;
        RECT 1478.870 1487.130 1481.770 1487.190 ;
        RECT 1658.870 1487.130 1661.770 1487.190 ;
        RECT 1838.870 1487.130 1841.770 1487.190 ;
        RECT 2018.870 1487.130 2021.770 1487.190 ;
        RECT 2198.870 1487.130 2201.770 1487.190 ;
        RECT 2378.870 1487.130 2381.770 1487.190 ;
        RECT 2558.870 1487.130 2561.770 1487.190 ;
        RECT 2738.870 1487.130 2741.770 1487.190 ;
        RECT 2945.050 1487.130 2947.950 1487.190 ;
        RECT -32.930 1484.230 2952.550 1487.130 ;
        RECT -28.330 1484.170 -25.430 1484.230 ;
        RECT 38.870 1484.170 41.770 1484.230 ;
        RECT 218.870 1484.170 221.770 1484.230 ;
        RECT 398.870 1484.170 401.770 1484.230 ;
        RECT 578.870 1484.170 581.770 1484.230 ;
        RECT 758.870 1484.170 761.770 1484.230 ;
        RECT 938.870 1484.170 941.770 1484.230 ;
        RECT 1118.870 1484.170 1121.770 1484.230 ;
        RECT 1298.870 1484.170 1301.770 1484.230 ;
        RECT 1478.870 1484.170 1481.770 1484.230 ;
        RECT 1658.870 1484.170 1661.770 1484.230 ;
        RECT 1838.870 1484.170 1841.770 1484.230 ;
        RECT 2018.870 1484.170 2021.770 1484.230 ;
        RECT 2198.870 1484.170 2201.770 1484.230 ;
        RECT 2378.870 1484.170 2381.770 1484.230 ;
        RECT 2558.870 1484.170 2561.770 1484.230 ;
        RECT 2738.870 1484.170 2741.770 1484.230 ;
        RECT 2945.050 1484.170 2947.950 1484.230 ;
        RECT -28.330 1307.130 -25.430 1307.190 ;
        RECT 38.870 1307.130 41.770 1307.190 ;
        RECT 218.870 1307.130 221.770 1307.190 ;
        RECT 398.870 1307.130 401.770 1307.190 ;
        RECT 578.870 1307.130 581.770 1307.190 ;
        RECT 758.870 1307.130 761.770 1307.190 ;
        RECT 938.870 1307.130 941.770 1307.190 ;
        RECT 1118.870 1307.130 1121.770 1307.190 ;
        RECT 1298.870 1307.130 1301.770 1307.190 ;
        RECT 1478.870 1307.130 1481.770 1307.190 ;
        RECT 1658.870 1307.130 1661.770 1307.190 ;
        RECT 1838.870 1307.130 1841.770 1307.190 ;
        RECT 2018.870 1307.130 2021.770 1307.190 ;
        RECT 2198.870 1307.130 2201.770 1307.190 ;
        RECT 2378.870 1307.130 2381.770 1307.190 ;
        RECT 2558.870 1307.130 2561.770 1307.190 ;
        RECT 2738.870 1307.130 2741.770 1307.190 ;
        RECT 2945.050 1307.130 2947.950 1307.190 ;
        RECT -32.930 1304.230 2952.550 1307.130 ;
        RECT -28.330 1304.170 -25.430 1304.230 ;
        RECT 38.870 1304.170 41.770 1304.230 ;
        RECT 218.870 1304.170 221.770 1304.230 ;
        RECT 398.870 1304.170 401.770 1304.230 ;
        RECT 578.870 1304.170 581.770 1304.230 ;
        RECT 758.870 1304.170 761.770 1304.230 ;
        RECT 938.870 1304.170 941.770 1304.230 ;
        RECT 1118.870 1304.170 1121.770 1304.230 ;
        RECT 1298.870 1304.170 1301.770 1304.230 ;
        RECT 1478.870 1304.170 1481.770 1304.230 ;
        RECT 1658.870 1304.170 1661.770 1304.230 ;
        RECT 1838.870 1304.170 1841.770 1304.230 ;
        RECT 2018.870 1304.170 2021.770 1304.230 ;
        RECT 2198.870 1304.170 2201.770 1304.230 ;
        RECT 2378.870 1304.170 2381.770 1304.230 ;
        RECT 2558.870 1304.170 2561.770 1304.230 ;
        RECT 2738.870 1304.170 2741.770 1304.230 ;
        RECT 2945.050 1304.170 2947.950 1304.230 ;
        RECT -28.330 1127.130 -25.430 1127.190 ;
        RECT 38.870 1127.130 41.770 1127.190 ;
        RECT 218.870 1127.130 221.770 1127.190 ;
        RECT 398.870 1127.130 401.770 1127.190 ;
        RECT 578.870 1127.130 581.770 1127.190 ;
        RECT 758.870 1127.130 761.770 1127.190 ;
        RECT 938.870 1127.130 941.770 1127.190 ;
        RECT 1118.870 1127.130 1121.770 1127.190 ;
        RECT 1298.870 1127.130 1301.770 1127.190 ;
        RECT 1478.870 1127.130 1481.770 1127.190 ;
        RECT 1658.870 1127.130 1661.770 1127.190 ;
        RECT 1838.870 1127.130 1841.770 1127.190 ;
        RECT 2018.870 1127.130 2021.770 1127.190 ;
        RECT 2198.870 1127.130 2201.770 1127.190 ;
        RECT 2378.870 1127.130 2381.770 1127.190 ;
        RECT 2558.870 1127.130 2561.770 1127.190 ;
        RECT 2738.870 1127.130 2741.770 1127.190 ;
        RECT 2945.050 1127.130 2947.950 1127.190 ;
        RECT -32.930 1124.230 2952.550 1127.130 ;
        RECT -28.330 1124.170 -25.430 1124.230 ;
        RECT 38.870 1124.170 41.770 1124.230 ;
        RECT 218.870 1124.170 221.770 1124.230 ;
        RECT 398.870 1124.170 401.770 1124.230 ;
        RECT 578.870 1124.170 581.770 1124.230 ;
        RECT 758.870 1124.170 761.770 1124.230 ;
        RECT 938.870 1124.170 941.770 1124.230 ;
        RECT 1118.870 1124.170 1121.770 1124.230 ;
        RECT 1298.870 1124.170 1301.770 1124.230 ;
        RECT 1478.870 1124.170 1481.770 1124.230 ;
        RECT 1658.870 1124.170 1661.770 1124.230 ;
        RECT 1838.870 1124.170 1841.770 1124.230 ;
        RECT 2018.870 1124.170 2021.770 1124.230 ;
        RECT 2198.870 1124.170 2201.770 1124.230 ;
        RECT 2378.870 1124.170 2381.770 1124.230 ;
        RECT 2558.870 1124.170 2561.770 1124.230 ;
        RECT 2738.870 1124.170 2741.770 1124.230 ;
        RECT 2945.050 1124.170 2947.950 1124.230 ;
        RECT -28.330 947.130 -25.430 947.190 ;
        RECT 38.870 947.130 41.770 947.190 ;
        RECT 218.870 947.130 221.770 947.190 ;
        RECT 398.870 947.130 401.770 947.190 ;
        RECT 578.870 947.130 581.770 947.190 ;
        RECT 758.870 947.130 761.770 947.190 ;
        RECT 938.870 947.130 941.770 947.190 ;
        RECT 1118.870 947.130 1121.770 947.190 ;
        RECT 1298.870 947.130 1301.770 947.190 ;
        RECT 1478.870 947.130 1481.770 947.190 ;
        RECT 1658.870 947.130 1661.770 947.190 ;
        RECT 1838.870 947.130 1841.770 947.190 ;
        RECT 2018.870 947.130 2021.770 947.190 ;
        RECT 2198.870 947.130 2201.770 947.190 ;
        RECT 2378.870 947.130 2381.770 947.190 ;
        RECT 2558.870 947.130 2561.770 947.190 ;
        RECT 2738.870 947.130 2741.770 947.190 ;
        RECT 2945.050 947.130 2947.950 947.190 ;
        RECT -32.930 944.230 2952.550 947.130 ;
        RECT -28.330 944.170 -25.430 944.230 ;
        RECT 38.870 944.170 41.770 944.230 ;
        RECT 218.870 944.170 221.770 944.230 ;
        RECT 398.870 944.170 401.770 944.230 ;
        RECT 578.870 944.170 581.770 944.230 ;
        RECT 758.870 944.170 761.770 944.230 ;
        RECT 938.870 944.170 941.770 944.230 ;
        RECT 1118.870 944.170 1121.770 944.230 ;
        RECT 1298.870 944.170 1301.770 944.230 ;
        RECT 1478.870 944.170 1481.770 944.230 ;
        RECT 1658.870 944.170 1661.770 944.230 ;
        RECT 1838.870 944.170 1841.770 944.230 ;
        RECT 2018.870 944.170 2021.770 944.230 ;
        RECT 2198.870 944.170 2201.770 944.230 ;
        RECT 2378.870 944.170 2381.770 944.230 ;
        RECT 2558.870 944.170 2561.770 944.230 ;
        RECT 2738.870 944.170 2741.770 944.230 ;
        RECT 2945.050 944.170 2947.950 944.230 ;
        RECT -28.330 767.130 -25.430 767.190 ;
        RECT 38.870 767.130 41.770 767.190 ;
        RECT 218.870 767.130 221.770 767.190 ;
        RECT 398.870 767.130 401.770 767.190 ;
        RECT 578.870 767.130 581.770 767.190 ;
        RECT 758.870 767.130 761.770 767.190 ;
        RECT 938.870 767.130 941.770 767.190 ;
        RECT 1118.870 767.130 1121.770 767.190 ;
        RECT 1298.870 767.130 1301.770 767.190 ;
        RECT 1478.870 767.130 1481.770 767.190 ;
        RECT 1658.870 767.130 1661.770 767.190 ;
        RECT 1838.870 767.130 1841.770 767.190 ;
        RECT 2018.870 767.130 2021.770 767.190 ;
        RECT 2198.870 767.130 2201.770 767.190 ;
        RECT 2378.870 767.130 2381.770 767.190 ;
        RECT 2558.870 767.130 2561.770 767.190 ;
        RECT 2738.870 767.130 2741.770 767.190 ;
        RECT 2945.050 767.130 2947.950 767.190 ;
        RECT -32.930 764.230 2952.550 767.130 ;
        RECT -28.330 764.170 -25.430 764.230 ;
        RECT 38.870 764.170 41.770 764.230 ;
        RECT 218.870 764.170 221.770 764.230 ;
        RECT 398.870 764.170 401.770 764.230 ;
        RECT 578.870 764.170 581.770 764.230 ;
        RECT 758.870 764.170 761.770 764.230 ;
        RECT 938.870 764.170 941.770 764.230 ;
        RECT 1118.870 764.170 1121.770 764.230 ;
        RECT 1298.870 764.170 1301.770 764.230 ;
        RECT 1478.870 764.170 1481.770 764.230 ;
        RECT 1658.870 764.170 1661.770 764.230 ;
        RECT 1838.870 764.170 1841.770 764.230 ;
        RECT 2018.870 764.170 2021.770 764.230 ;
        RECT 2198.870 764.170 2201.770 764.230 ;
        RECT 2378.870 764.170 2381.770 764.230 ;
        RECT 2558.870 764.170 2561.770 764.230 ;
        RECT 2738.870 764.170 2741.770 764.230 ;
        RECT 2945.050 764.170 2947.950 764.230 ;
        RECT -28.330 587.130 -25.430 587.190 ;
        RECT 38.870 587.130 41.770 587.190 ;
        RECT 218.870 587.130 221.770 587.190 ;
        RECT 398.870 587.130 401.770 587.190 ;
        RECT 578.870 587.130 581.770 587.190 ;
        RECT 758.870 587.130 761.770 587.190 ;
        RECT 938.870 587.130 941.770 587.190 ;
        RECT 1118.870 587.130 1121.770 587.190 ;
        RECT 1298.870 587.130 1301.770 587.190 ;
        RECT 1478.870 587.130 1481.770 587.190 ;
        RECT 1658.870 587.130 1661.770 587.190 ;
        RECT 1838.870 587.130 1841.770 587.190 ;
        RECT 2018.870 587.130 2021.770 587.190 ;
        RECT 2198.870 587.130 2201.770 587.190 ;
        RECT 2378.870 587.130 2381.770 587.190 ;
        RECT 2558.870 587.130 2561.770 587.190 ;
        RECT 2738.870 587.130 2741.770 587.190 ;
        RECT 2945.050 587.130 2947.950 587.190 ;
        RECT -32.930 584.230 2952.550 587.130 ;
        RECT -28.330 584.170 -25.430 584.230 ;
        RECT 38.870 584.170 41.770 584.230 ;
        RECT 218.870 584.170 221.770 584.230 ;
        RECT 398.870 584.170 401.770 584.230 ;
        RECT 578.870 584.170 581.770 584.230 ;
        RECT 758.870 584.170 761.770 584.230 ;
        RECT 938.870 584.170 941.770 584.230 ;
        RECT 1118.870 584.170 1121.770 584.230 ;
        RECT 1298.870 584.170 1301.770 584.230 ;
        RECT 1478.870 584.170 1481.770 584.230 ;
        RECT 1658.870 584.170 1661.770 584.230 ;
        RECT 1838.870 584.170 1841.770 584.230 ;
        RECT 2018.870 584.170 2021.770 584.230 ;
        RECT 2198.870 584.170 2201.770 584.230 ;
        RECT 2378.870 584.170 2381.770 584.230 ;
        RECT 2558.870 584.170 2561.770 584.230 ;
        RECT 2738.870 584.170 2741.770 584.230 ;
        RECT 2945.050 584.170 2947.950 584.230 ;
        RECT -28.330 407.130 -25.430 407.190 ;
        RECT 38.870 407.130 41.770 407.190 ;
        RECT 218.870 407.130 221.770 407.190 ;
        RECT 398.870 407.130 401.770 407.190 ;
        RECT 578.870 407.130 581.770 407.190 ;
        RECT 758.870 407.130 761.770 407.190 ;
        RECT 938.870 407.130 941.770 407.190 ;
        RECT 1118.870 407.130 1121.770 407.190 ;
        RECT 1298.870 407.130 1301.770 407.190 ;
        RECT 1478.870 407.130 1481.770 407.190 ;
        RECT 1658.870 407.130 1661.770 407.190 ;
        RECT 1838.870 407.130 1841.770 407.190 ;
        RECT 2018.870 407.130 2021.770 407.190 ;
        RECT 2198.870 407.130 2201.770 407.190 ;
        RECT 2378.870 407.130 2381.770 407.190 ;
        RECT 2558.870 407.130 2561.770 407.190 ;
        RECT 2738.870 407.130 2741.770 407.190 ;
        RECT 2945.050 407.130 2947.950 407.190 ;
        RECT -32.930 404.230 2952.550 407.130 ;
        RECT -28.330 404.170 -25.430 404.230 ;
        RECT 38.870 404.170 41.770 404.230 ;
        RECT 218.870 404.170 221.770 404.230 ;
        RECT 398.870 404.170 401.770 404.230 ;
        RECT 578.870 404.170 581.770 404.230 ;
        RECT 758.870 404.170 761.770 404.230 ;
        RECT 938.870 404.170 941.770 404.230 ;
        RECT 1118.870 404.170 1121.770 404.230 ;
        RECT 1298.870 404.170 1301.770 404.230 ;
        RECT 1478.870 404.170 1481.770 404.230 ;
        RECT 1658.870 404.170 1661.770 404.230 ;
        RECT 1838.870 404.170 1841.770 404.230 ;
        RECT 2018.870 404.170 2021.770 404.230 ;
        RECT 2198.870 404.170 2201.770 404.230 ;
        RECT 2378.870 404.170 2381.770 404.230 ;
        RECT 2558.870 404.170 2561.770 404.230 ;
        RECT 2738.870 404.170 2741.770 404.230 ;
        RECT 2945.050 404.170 2947.950 404.230 ;
        RECT -28.330 227.130 -25.430 227.190 ;
        RECT 38.870 227.130 41.770 227.190 ;
        RECT 218.870 227.130 221.770 227.190 ;
        RECT 398.870 227.130 401.770 227.190 ;
        RECT 578.870 227.130 581.770 227.190 ;
        RECT 758.870 227.130 761.770 227.190 ;
        RECT 938.870 227.130 941.770 227.190 ;
        RECT 1118.870 227.130 1121.770 227.190 ;
        RECT 1298.870 227.130 1301.770 227.190 ;
        RECT 1478.870 227.130 1481.770 227.190 ;
        RECT 1658.870 227.130 1661.770 227.190 ;
        RECT 1838.870 227.130 1841.770 227.190 ;
        RECT 2018.870 227.130 2021.770 227.190 ;
        RECT 2198.870 227.130 2201.770 227.190 ;
        RECT 2378.870 227.130 2381.770 227.190 ;
        RECT 2558.870 227.130 2561.770 227.190 ;
        RECT 2738.870 227.130 2741.770 227.190 ;
        RECT 2945.050 227.130 2947.950 227.190 ;
        RECT -32.930 224.230 2952.550 227.130 ;
        RECT -28.330 224.170 -25.430 224.230 ;
        RECT 38.870 224.170 41.770 224.230 ;
        RECT 218.870 224.170 221.770 224.230 ;
        RECT 398.870 224.170 401.770 224.230 ;
        RECT 578.870 224.170 581.770 224.230 ;
        RECT 758.870 224.170 761.770 224.230 ;
        RECT 938.870 224.170 941.770 224.230 ;
        RECT 1118.870 224.170 1121.770 224.230 ;
        RECT 1298.870 224.170 1301.770 224.230 ;
        RECT 1478.870 224.170 1481.770 224.230 ;
        RECT 1658.870 224.170 1661.770 224.230 ;
        RECT 1838.870 224.170 1841.770 224.230 ;
        RECT 2018.870 224.170 2021.770 224.230 ;
        RECT 2198.870 224.170 2201.770 224.230 ;
        RECT 2378.870 224.170 2381.770 224.230 ;
        RECT 2558.870 224.170 2561.770 224.230 ;
        RECT 2738.870 224.170 2741.770 224.230 ;
        RECT 2945.050 224.170 2947.950 224.230 ;
        RECT -28.330 47.130 -25.430 47.190 ;
        RECT 38.870 47.130 41.770 47.190 ;
        RECT 218.870 47.130 221.770 47.190 ;
        RECT 398.870 47.130 401.770 47.190 ;
        RECT 578.870 47.130 581.770 47.190 ;
        RECT 758.870 47.130 761.770 47.190 ;
        RECT 938.870 47.130 941.770 47.190 ;
        RECT 1118.870 47.130 1121.770 47.190 ;
        RECT 1298.870 47.130 1301.770 47.190 ;
        RECT 1478.870 47.130 1481.770 47.190 ;
        RECT 1658.870 47.130 1661.770 47.190 ;
        RECT 1838.870 47.130 1841.770 47.190 ;
        RECT 2018.870 47.130 2021.770 47.190 ;
        RECT 2198.870 47.130 2201.770 47.190 ;
        RECT 2378.870 47.130 2381.770 47.190 ;
        RECT 2558.870 47.130 2561.770 47.190 ;
        RECT 2738.870 47.130 2741.770 47.190 ;
        RECT 2945.050 47.130 2947.950 47.190 ;
        RECT -32.930 44.230 2952.550 47.130 ;
        RECT -28.330 44.170 -25.430 44.230 ;
        RECT 38.870 44.170 41.770 44.230 ;
        RECT 218.870 44.170 221.770 44.230 ;
        RECT 398.870 44.170 401.770 44.230 ;
        RECT 578.870 44.170 581.770 44.230 ;
        RECT 758.870 44.170 761.770 44.230 ;
        RECT 938.870 44.170 941.770 44.230 ;
        RECT 1118.870 44.170 1121.770 44.230 ;
        RECT 1298.870 44.170 1301.770 44.230 ;
        RECT 1478.870 44.170 1481.770 44.230 ;
        RECT 1658.870 44.170 1661.770 44.230 ;
        RECT 1838.870 44.170 1841.770 44.230 ;
        RECT 2018.870 44.170 2021.770 44.230 ;
        RECT 2198.870 44.170 2201.770 44.230 ;
        RECT 2378.870 44.170 2381.770 44.230 ;
        RECT 2558.870 44.170 2561.770 44.230 ;
        RECT 2738.870 44.170 2741.770 44.230 ;
        RECT 2945.050 44.170 2947.950 44.230 ;
        RECT -28.330 -20.070 -25.430 -20.010 ;
        RECT 38.870 -20.070 41.770 -20.010 ;
        RECT 218.870 -20.070 221.770 -20.010 ;
        RECT 398.870 -20.070 401.770 -20.010 ;
        RECT 578.870 -20.070 581.770 -20.010 ;
        RECT 758.870 -20.070 761.770 -20.010 ;
        RECT 938.870 -20.070 941.770 -20.010 ;
        RECT 1118.870 -20.070 1121.770 -20.010 ;
        RECT 1298.870 -20.070 1301.770 -20.010 ;
        RECT 1478.870 -20.070 1481.770 -20.010 ;
        RECT 1658.870 -20.070 1661.770 -20.010 ;
        RECT 1838.870 -20.070 1841.770 -20.010 ;
        RECT 2018.870 -20.070 2021.770 -20.010 ;
        RECT 2198.870 -20.070 2201.770 -20.010 ;
        RECT 2378.870 -20.070 2381.770 -20.010 ;
        RECT 2558.870 -20.070 2561.770 -20.010 ;
        RECT 2738.870 -20.070 2741.770 -20.010 ;
        RECT 2945.050 -20.070 2947.950 -20.010 ;
        RECT -28.330 -22.970 2947.950 -20.070 ;
        RECT -28.330 -23.030 -25.430 -22.970 ;
        RECT 38.870 -23.030 41.770 -22.970 ;
        RECT 218.870 -23.030 221.770 -22.970 ;
        RECT 398.870 -23.030 401.770 -22.970 ;
        RECT 578.870 -23.030 581.770 -22.970 ;
        RECT 758.870 -23.030 761.770 -22.970 ;
        RECT 938.870 -23.030 941.770 -22.970 ;
        RECT 1118.870 -23.030 1121.770 -22.970 ;
        RECT 1298.870 -23.030 1301.770 -22.970 ;
        RECT 1478.870 -23.030 1481.770 -22.970 ;
        RECT 1658.870 -23.030 1661.770 -22.970 ;
        RECT 1838.870 -23.030 1841.770 -22.970 ;
        RECT 2018.870 -23.030 2021.770 -22.970 ;
        RECT 2198.870 -23.030 2201.770 -22.970 ;
        RECT 2378.870 -23.030 2381.770 -22.970 ;
        RECT 2558.870 -23.030 2561.770 -22.970 ;
        RECT 2738.870 -23.030 2741.770 -22.970 ;
        RECT 2945.050 -23.030 2947.950 -22.970 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.930 -27.570 -30.030 3547.250 ;
        RECT 128.870 -27.570 131.770 3547.250 ;
        RECT 308.870 -27.570 311.770 3547.250 ;
        RECT 488.870 -27.570 491.770 3547.250 ;
        RECT 668.870 -27.570 671.770 3547.250 ;
        RECT 848.870 -27.570 851.770 3547.250 ;
        RECT 1028.870 -27.570 1031.770 3547.250 ;
        RECT 1208.870 -27.570 1211.770 3547.250 ;
        RECT 1388.870 -27.570 1391.770 3547.250 ;
        RECT 1568.870 -27.570 1571.770 3547.250 ;
        RECT 1748.870 -27.570 1751.770 3547.250 ;
        RECT 1928.870 -27.570 1931.770 3547.250 ;
        RECT 2108.870 -27.570 2111.770 3547.250 ;
        RECT 2288.870 -27.570 2291.770 3547.250 ;
        RECT 2468.870 -27.570 2471.770 3547.250 ;
        RECT 2648.870 -27.570 2651.770 3547.250 ;
        RECT 2828.870 -27.570 2831.770 3547.250 ;
        RECT 2949.650 -27.570 2952.550 3547.250 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3375.890 -30.890 3377.070 ;
        RECT -32.070 3374.290 -30.890 3375.470 ;
        RECT -32.070 3195.890 -30.890 3197.070 ;
        RECT -32.070 3194.290 -30.890 3195.470 ;
        RECT -32.070 3015.890 -30.890 3017.070 ;
        RECT -32.070 3014.290 -30.890 3015.470 ;
        RECT -32.070 2835.890 -30.890 2837.070 ;
        RECT -32.070 2834.290 -30.890 2835.470 ;
        RECT -32.070 2655.890 -30.890 2657.070 ;
        RECT -32.070 2654.290 -30.890 2655.470 ;
        RECT -32.070 2475.890 -30.890 2477.070 ;
        RECT -32.070 2474.290 -30.890 2475.470 ;
        RECT -32.070 2295.890 -30.890 2297.070 ;
        RECT -32.070 2294.290 -30.890 2295.470 ;
        RECT -32.070 2115.890 -30.890 2117.070 ;
        RECT -32.070 2114.290 -30.890 2115.470 ;
        RECT -32.070 1935.890 -30.890 1937.070 ;
        RECT -32.070 1934.290 -30.890 1935.470 ;
        RECT -32.070 1755.890 -30.890 1757.070 ;
        RECT -32.070 1754.290 -30.890 1755.470 ;
        RECT -32.070 1575.890 -30.890 1577.070 ;
        RECT -32.070 1574.290 -30.890 1575.470 ;
        RECT -32.070 1395.890 -30.890 1397.070 ;
        RECT -32.070 1394.290 -30.890 1395.470 ;
        RECT -32.070 1215.890 -30.890 1217.070 ;
        RECT -32.070 1214.290 -30.890 1215.470 ;
        RECT -32.070 1035.890 -30.890 1037.070 ;
        RECT -32.070 1034.290 -30.890 1035.470 ;
        RECT -32.070 855.890 -30.890 857.070 ;
        RECT -32.070 854.290 -30.890 855.470 ;
        RECT -32.070 675.890 -30.890 677.070 ;
        RECT -32.070 674.290 -30.890 675.470 ;
        RECT -32.070 495.890 -30.890 497.070 ;
        RECT -32.070 494.290 -30.890 495.470 ;
        RECT -32.070 315.890 -30.890 317.070 ;
        RECT -32.070 314.290 -30.890 315.470 ;
        RECT -32.070 135.890 -30.890 137.070 ;
        RECT -32.070 134.290 -30.890 135.470 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 129.730 3546.010 130.910 3547.190 ;
        RECT 129.730 3544.410 130.910 3545.590 ;
        RECT 129.730 3375.890 130.910 3377.070 ;
        RECT 129.730 3374.290 130.910 3375.470 ;
        RECT 129.730 3195.890 130.910 3197.070 ;
        RECT 129.730 3194.290 130.910 3195.470 ;
        RECT 129.730 3015.890 130.910 3017.070 ;
        RECT 129.730 3014.290 130.910 3015.470 ;
        RECT 129.730 2835.890 130.910 2837.070 ;
        RECT 129.730 2834.290 130.910 2835.470 ;
        RECT 129.730 2655.890 130.910 2657.070 ;
        RECT 129.730 2654.290 130.910 2655.470 ;
        RECT 129.730 2475.890 130.910 2477.070 ;
        RECT 129.730 2474.290 130.910 2475.470 ;
        RECT 129.730 2295.890 130.910 2297.070 ;
        RECT 129.730 2294.290 130.910 2295.470 ;
        RECT 129.730 2115.890 130.910 2117.070 ;
        RECT 129.730 2114.290 130.910 2115.470 ;
        RECT 129.730 1935.890 130.910 1937.070 ;
        RECT 129.730 1934.290 130.910 1935.470 ;
        RECT 129.730 1755.890 130.910 1757.070 ;
        RECT 129.730 1754.290 130.910 1755.470 ;
        RECT 129.730 1575.890 130.910 1577.070 ;
        RECT 129.730 1574.290 130.910 1575.470 ;
        RECT 129.730 1395.890 130.910 1397.070 ;
        RECT 129.730 1394.290 130.910 1395.470 ;
        RECT 129.730 1215.890 130.910 1217.070 ;
        RECT 129.730 1214.290 130.910 1215.470 ;
        RECT 129.730 1035.890 130.910 1037.070 ;
        RECT 129.730 1034.290 130.910 1035.470 ;
        RECT 129.730 855.890 130.910 857.070 ;
        RECT 129.730 854.290 130.910 855.470 ;
        RECT 129.730 675.890 130.910 677.070 ;
        RECT 129.730 674.290 130.910 675.470 ;
        RECT 129.730 495.890 130.910 497.070 ;
        RECT 129.730 494.290 130.910 495.470 ;
        RECT 129.730 315.890 130.910 317.070 ;
        RECT 129.730 314.290 130.910 315.470 ;
        RECT 129.730 135.890 130.910 137.070 ;
        RECT 129.730 134.290 130.910 135.470 ;
        RECT 129.730 -25.910 130.910 -24.730 ;
        RECT 129.730 -27.510 130.910 -26.330 ;
        RECT 309.730 3546.010 310.910 3547.190 ;
        RECT 309.730 3544.410 310.910 3545.590 ;
        RECT 309.730 3375.890 310.910 3377.070 ;
        RECT 309.730 3374.290 310.910 3375.470 ;
        RECT 309.730 3195.890 310.910 3197.070 ;
        RECT 309.730 3194.290 310.910 3195.470 ;
        RECT 309.730 3015.890 310.910 3017.070 ;
        RECT 309.730 3014.290 310.910 3015.470 ;
        RECT 309.730 2835.890 310.910 2837.070 ;
        RECT 309.730 2834.290 310.910 2835.470 ;
        RECT 309.730 2655.890 310.910 2657.070 ;
        RECT 309.730 2654.290 310.910 2655.470 ;
        RECT 309.730 2475.890 310.910 2477.070 ;
        RECT 309.730 2474.290 310.910 2475.470 ;
        RECT 309.730 2295.890 310.910 2297.070 ;
        RECT 309.730 2294.290 310.910 2295.470 ;
        RECT 309.730 2115.890 310.910 2117.070 ;
        RECT 309.730 2114.290 310.910 2115.470 ;
        RECT 309.730 1935.890 310.910 1937.070 ;
        RECT 309.730 1934.290 310.910 1935.470 ;
        RECT 309.730 1755.890 310.910 1757.070 ;
        RECT 309.730 1754.290 310.910 1755.470 ;
        RECT 309.730 1575.890 310.910 1577.070 ;
        RECT 309.730 1574.290 310.910 1575.470 ;
        RECT 309.730 1395.890 310.910 1397.070 ;
        RECT 309.730 1394.290 310.910 1395.470 ;
        RECT 309.730 1215.890 310.910 1217.070 ;
        RECT 309.730 1214.290 310.910 1215.470 ;
        RECT 309.730 1035.890 310.910 1037.070 ;
        RECT 309.730 1034.290 310.910 1035.470 ;
        RECT 309.730 855.890 310.910 857.070 ;
        RECT 309.730 854.290 310.910 855.470 ;
        RECT 309.730 675.890 310.910 677.070 ;
        RECT 309.730 674.290 310.910 675.470 ;
        RECT 309.730 495.890 310.910 497.070 ;
        RECT 309.730 494.290 310.910 495.470 ;
        RECT 309.730 315.890 310.910 317.070 ;
        RECT 309.730 314.290 310.910 315.470 ;
        RECT 309.730 135.890 310.910 137.070 ;
        RECT 309.730 134.290 310.910 135.470 ;
        RECT 309.730 -25.910 310.910 -24.730 ;
        RECT 309.730 -27.510 310.910 -26.330 ;
        RECT 489.730 3546.010 490.910 3547.190 ;
        RECT 489.730 3544.410 490.910 3545.590 ;
        RECT 489.730 3375.890 490.910 3377.070 ;
        RECT 489.730 3374.290 490.910 3375.470 ;
        RECT 489.730 3195.890 490.910 3197.070 ;
        RECT 489.730 3194.290 490.910 3195.470 ;
        RECT 489.730 3015.890 490.910 3017.070 ;
        RECT 489.730 3014.290 490.910 3015.470 ;
        RECT 489.730 2835.890 490.910 2837.070 ;
        RECT 489.730 2834.290 490.910 2835.470 ;
        RECT 489.730 2655.890 490.910 2657.070 ;
        RECT 489.730 2654.290 490.910 2655.470 ;
        RECT 489.730 2475.890 490.910 2477.070 ;
        RECT 489.730 2474.290 490.910 2475.470 ;
        RECT 489.730 2295.890 490.910 2297.070 ;
        RECT 489.730 2294.290 490.910 2295.470 ;
        RECT 489.730 2115.890 490.910 2117.070 ;
        RECT 489.730 2114.290 490.910 2115.470 ;
        RECT 489.730 1935.890 490.910 1937.070 ;
        RECT 489.730 1934.290 490.910 1935.470 ;
        RECT 489.730 1755.890 490.910 1757.070 ;
        RECT 489.730 1754.290 490.910 1755.470 ;
        RECT 489.730 1575.890 490.910 1577.070 ;
        RECT 489.730 1574.290 490.910 1575.470 ;
        RECT 489.730 1395.890 490.910 1397.070 ;
        RECT 489.730 1394.290 490.910 1395.470 ;
        RECT 489.730 1215.890 490.910 1217.070 ;
        RECT 489.730 1214.290 490.910 1215.470 ;
        RECT 489.730 1035.890 490.910 1037.070 ;
        RECT 489.730 1034.290 490.910 1035.470 ;
        RECT 489.730 855.890 490.910 857.070 ;
        RECT 489.730 854.290 490.910 855.470 ;
        RECT 489.730 675.890 490.910 677.070 ;
        RECT 489.730 674.290 490.910 675.470 ;
        RECT 489.730 495.890 490.910 497.070 ;
        RECT 489.730 494.290 490.910 495.470 ;
        RECT 489.730 315.890 490.910 317.070 ;
        RECT 489.730 314.290 490.910 315.470 ;
        RECT 489.730 135.890 490.910 137.070 ;
        RECT 489.730 134.290 490.910 135.470 ;
        RECT 489.730 -25.910 490.910 -24.730 ;
        RECT 489.730 -27.510 490.910 -26.330 ;
        RECT 669.730 3546.010 670.910 3547.190 ;
        RECT 669.730 3544.410 670.910 3545.590 ;
        RECT 669.730 3375.890 670.910 3377.070 ;
        RECT 669.730 3374.290 670.910 3375.470 ;
        RECT 669.730 3195.890 670.910 3197.070 ;
        RECT 669.730 3194.290 670.910 3195.470 ;
        RECT 669.730 3015.890 670.910 3017.070 ;
        RECT 669.730 3014.290 670.910 3015.470 ;
        RECT 669.730 2835.890 670.910 2837.070 ;
        RECT 669.730 2834.290 670.910 2835.470 ;
        RECT 669.730 2655.890 670.910 2657.070 ;
        RECT 669.730 2654.290 670.910 2655.470 ;
        RECT 669.730 2475.890 670.910 2477.070 ;
        RECT 669.730 2474.290 670.910 2475.470 ;
        RECT 669.730 2295.890 670.910 2297.070 ;
        RECT 669.730 2294.290 670.910 2295.470 ;
        RECT 669.730 2115.890 670.910 2117.070 ;
        RECT 669.730 2114.290 670.910 2115.470 ;
        RECT 669.730 1935.890 670.910 1937.070 ;
        RECT 669.730 1934.290 670.910 1935.470 ;
        RECT 669.730 1755.890 670.910 1757.070 ;
        RECT 669.730 1754.290 670.910 1755.470 ;
        RECT 669.730 1575.890 670.910 1577.070 ;
        RECT 669.730 1574.290 670.910 1575.470 ;
        RECT 669.730 1395.890 670.910 1397.070 ;
        RECT 669.730 1394.290 670.910 1395.470 ;
        RECT 669.730 1215.890 670.910 1217.070 ;
        RECT 669.730 1214.290 670.910 1215.470 ;
        RECT 669.730 1035.890 670.910 1037.070 ;
        RECT 669.730 1034.290 670.910 1035.470 ;
        RECT 669.730 855.890 670.910 857.070 ;
        RECT 669.730 854.290 670.910 855.470 ;
        RECT 669.730 675.890 670.910 677.070 ;
        RECT 669.730 674.290 670.910 675.470 ;
        RECT 669.730 495.890 670.910 497.070 ;
        RECT 669.730 494.290 670.910 495.470 ;
        RECT 669.730 315.890 670.910 317.070 ;
        RECT 669.730 314.290 670.910 315.470 ;
        RECT 669.730 135.890 670.910 137.070 ;
        RECT 669.730 134.290 670.910 135.470 ;
        RECT 669.730 -25.910 670.910 -24.730 ;
        RECT 669.730 -27.510 670.910 -26.330 ;
        RECT 849.730 3546.010 850.910 3547.190 ;
        RECT 849.730 3544.410 850.910 3545.590 ;
        RECT 849.730 3375.890 850.910 3377.070 ;
        RECT 849.730 3374.290 850.910 3375.470 ;
        RECT 849.730 3195.890 850.910 3197.070 ;
        RECT 849.730 3194.290 850.910 3195.470 ;
        RECT 849.730 3015.890 850.910 3017.070 ;
        RECT 849.730 3014.290 850.910 3015.470 ;
        RECT 849.730 2835.890 850.910 2837.070 ;
        RECT 849.730 2834.290 850.910 2835.470 ;
        RECT 849.730 2655.890 850.910 2657.070 ;
        RECT 849.730 2654.290 850.910 2655.470 ;
        RECT 849.730 2475.890 850.910 2477.070 ;
        RECT 849.730 2474.290 850.910 2475.470 ;
        RECT 849.730 2295.890 850.910 2297.070 ;
        RECT 849.730 2294.290 850.910 2295.470 ;
        RECT 849.730 2115.890 850.910 2117.070 ;
        RECT 849.730 2114.290 850.910 2115.470 ;
        RECT 849.730 1935.890 850.910 1937.070 ;
        RECT 849.730 1934.290 850.910 1935.470 ;
        RECT 849.730 1755.890 850.910 1757.070 ;
        RECT 849.730 1754.290 850.910 1755.470 ;
        RECT 849.730 1575.890 850.910 1577.070 ;
        RECT 849.730 1574.290 850.910 1575.470 ;
        RECT 849.730 1395.890 850.910 1397.070 ;
        RECT 849.730 1394.290 850.910 1395.470 ;
        RECT 849.730 1215.890 850.910 1217.070 ;
        RECT 849.730 1214.290 850.910 1215.470 ;
        RECT 849.730 1035.890 850.910 1037.070 ;
        RECT 849.730 1034.290 850.910 1035.470 ;
        RECT 849.730 855.890 850.910 857.070 ;
        RECT 849.730 854.290 850.910 855.470 ;
        RECT 849.730 675.890 850.910 677.070 ;
        RECT 849.730 674.290 850.910 675.470 ;
        RECT 849.730 495.890 850.910 497.070 ;
        RECT 849.730 494.290 850.910 495.470 ;
        RECT 849.730 315.890 850.910 317.070 ;
        RECT 849.730 314.290 850.910 315.470 ;
        RECT 849.730 135.890 850.910 137.070 ;
        RECT 849.730 134.290 850.910 135.470 ;
        RECT 849.730 -25.910 850.910 -24.730 ;
        RECT 849.730 -27.510 850.910 -26.330 ;
        RECT 1029.730 3546.010 1030.910 3547.190 ;
        RECT 1029.730 3544.410 1030.910 3545.590 ;
        RECT 1029.730 3375.890 1030.910 3377.070 ;
        RECT 1029.730 3374.290 1030.910 3375.470 ;
        RECT 1029.730 3195.890 1030.910 3197.070 ;
        RECT 1029.730 3194.290 1030.910 3195.470 ;
        RECT 1029.730 3015.890 1030.910 3017.070 ;
        RECT 1029.730 3014.290 1030.910 3015.470 ;
        RECT 1029.730 2835.890 1030.910 2837.070 ;
        RECT 1029.730 2834.290 1030.910 2835.470 ;
        RECT 1029.730 2655.890 1030.910 2657.070 ;
        RECT 1029.730 2654.290 1030.910 2655.470 ;
        RECT 1029.730 2475.890 1030.910 2477.070 ;
        RECT 1029.730 2474.290 1030.910 2475.470 ;
        RECT 1029.730 2295.890 1030.910 2297.070 ;
        RECT 1029.730 2294.290 1030.910 2295.470 ;
        RECT 1029.730 2115.890 1030.910 2117.070 ;
        RECT 1029.730 2114.290 1030.910 2115.470 ;
        RECT 1029.730 1935.890 1030.910 1937.070 ;
        RECT 1029.730 1934.290 1030.910 1935.470 ;
        RECT 1029.730 1755.890 1030.910 1757.070 ;
        RECT 1029.730 1754.290 1030.910 1755.470 ;
        RECT 1029.730 1575.890 1030.910 1577.070 ;
        RECT 1029.730 1574.290 1030.910 1575.470 ;
        RECT 1029.730 1395.890 1030.910 1397.070 ;
        RECT 1029.730 1394.290 1030.910 1395.470 ;
        RECT 1029.730 1215.890 1030.910 1217.070 ;
        RECT 1029.730 1214.290 1030.910 1215.470 ;
        RECT 1029.730 1035.890 1030.910 1037.070 ;
        RECT 1029.730 1034.290 1030.910 1035.470 ;
        RECT 1029.730 855.890 1030.910 857.070 ;
        RECT 1029.730 854.290 1030.910 855.470 ;
        RECT 1029.730 675.890 1030.910 677.070 ;
        RECT 1029.730 674.290 1030.910 675.470 ;
        RECT 1029.730 495.890 1030.910 497.070 ;
        RECT 1029.730 494.290 1030.910 495.470 ;
        RECT 1029.730 315.890 1030.910 317.070 ;
        RECT 1029.730 314.290 1030.910 315.470 ;
        RECT 1029.730 135.890 1030.910 137.070 ;
        RECT 1029.730 134.290 1030.910 135.470 ;
        RECT 1029.730 -25.910 1030.910 -24.730 ;
        RECT 1029.730 -27.510 1030.910 -26.330 ;
        RECT 1209.730 3546.010 1210.910 3547.190 ;
        RECT 1209.730 3544.410 1210.910 3545.590 ;
        RECT 1209.730 3375.890 1210.910 3377.070 ;
        RECT 1209.730 3374.290 1210.910 3375.470 ;
        RECT 1209.730 3195.890 1210.910 3197.070 ;
        RECT 1209.730 3194.290 1210.910 3195.470 ;
        RECT 1209.730 3015.890 1210.910 3017.070 ;
        RECT 1209.730 3014.290 1210.910 3015.470 ;
        RECT 1209.730 2835.890 1210.910 2837.070 ;
        RECT 1209.730 2834.290 1210.910 2835.470 ;
        RECT 1209.730 2655.890 1210.910 2657.070 ;
        RECT 1209.730 2654.290 1210.910 2655.470 ;
        RECT 1209.730 2475.890 1210.910 2477.070 ;
        RECT 1209.730 2474.290 1210.910 2475.470 ;
        RECT 1209.730 2295.890 1210.910 2297.070 ;
        RECT 1209.730 2294.290 1210.910 2295.470 ;
        RECT 1209.730 2115.890 1210.910 2117.070 ;
        RECT 1209.730 2114.290 1210.910 2115.470 ;
        RECT 1209.730 1935.890 1210.910 1937.070 ;
        RECT 1209.730 1934.290 1210.910 1935.470 ;
        RECT 1209.730 1755.890 1210.910 1757.070 ;
        RECT 1209.730 1754.290 1210.910 1755.470 ;
        RECT 1209.730 1575.890 1210.910 1577.070 ;
        RECT 1209.730 1574.290 1210.910 1575.470 ;
        RECT 1209.730 1395.890 1210.910 1397.070 ;
        RECT 1209.730 1394.290 1210.910 1395.470 ;
        RECT 1209.730 1215.890 1210.910 1217.070 ;
        RECT 1209.730 1214.290 1210.910 1215.470 ;
        RECT 1209.730 1035.890 1210.910 1037.070 ;
        RECT 1209.730 1034.290 1210.910 1035.470 ;
        RECT 1209.730 855.890 1210.910 857.070 ;
        RECT 1209.730 854.290 1210.910 855.470 ;
        RECT 1209.730 675.890 1210.910 677.070 ;
        RECT 1209.730 674.290 1210.910 675.470 ;
        RECT 1209.730 495.890 1210.910 497.070 ;
        RECT 1209.730 494.290 1210.910 495.470 ;
        RECT 1209.730 315.890 1210.910 317.070 ;
        RECT 1209.730 314.290 1210.910 315.470 ;
        RECT 1209.730 135.890 1210.910 137.070 ;
        RECT 1209.730 134.290 1210.910 135.470 ;
        RECT 1209.730 -25.910 1210.910 -24.730 ;
        RECT 1209.730 -27.510 1210.910 -26.330 ;
        RECT 1389.730 3546.010 1390.910 3547.190 ;
        RECT 1389.730 3544.410 1390.910 3545.590 ;
        RECT 1389.730 3375.890 1390.910 3377.070 ;
        RECT 1389.730 3374.290 1390.910 3375.470 ;
        RECT 1389.730 3195.890 1390.910 3197.070 ;
        RECT 1389.730 3194.290 1390.910 3195.470 ;
        RECT 1389.730 3015.890 1390.910 3017.070 ;
        RECT 1389.730 3014.290 1390.910 3015.470 ;
        RECT 1389.730 2835.890 1390.910 2837.070 ;
        RECT 1389.730 2834.290 1390.910 2835.470 ;
        RECT 1389.730 2655.890 1390.910 2657.070 ;
        RECT 1389.730 2654.290 1390.910 2655.470 ;
        RECT 1389.730 2475.890 1390.910 2477.070 ;
        RECT 1389.730 2474.290 1390.910 2475.470 ;
        RECT 1389.730 2295.890 1390.910 2297.070 ;
        RECT 1389.730 2294.290 1390.910 2295.470 ;
        RECT 1389.730 2115.890 1390.910 2117.070 ;
        RECT 1389.730 2114.290 1390.910 2115.470 ;
        RECT 1389.730 1935.890 1390.910 1937.070 ;
        RECT 1389.730 1934.290 1390.910 1935.470 ;
        RECT 1389.730 1755.890 1390.910 1757.070 ;
        RECT 1389.730 1754.290 1390.910 1755.470 ;
        RECT 1389.730 1575.890 1390.910 1577.070 ;
        RECT 1389.730 1574.290 1390.910 1575.470 ;
        RECT 1389.730 1395.890 1390.910 1397.070 ;
        RECT 1389.730 1394.290 1390.910 1395.470 ;
        RECT 1389.730 1215.890 1390.910 1217.070 ;
        RECT 1389.730 1214.290 1390.910 1215.470 ;
        RECT 1389.730 1035.890 1390.910 1037.070 ;
        RECT 1389.730 1034.290 1390.910 1035.470 ;
        RECT 1389.730 855.890 1390.910 857.070 ;
        RECT 1389.730 854.290 1390.910 855.470 ;
        RECT 1389.730 675.890 1390.910 677.070 ;
        RECT 1389.730 674.290 1390.910 675.470 ;
        RECT 1389.730 495.890 1390.910 497.070 ;
        RECT 1389.730 494.290 1390.910 495.470 ;
        RECT 1389.730 315.890 1390.910 317.070 ;
        RECT 1389.730 314.290 1390.910 315.470 ;
        RECT 1389.730 135.890 1390.910 137.070 ;
        RECT 1389.730 134.290 1390.910 135.470 ;
        RECT 1389.730 -25.910 1390.910 -24.730 ;
        RECT 1389.730 -27.510 1390.910 -26.330 ;
        RECT 1569.730 3546.010 1570.910 3547.190 ;
        RECT 1569.730 3544.410 1570.910 3545.590 ;
        RECT 1569.730 3375.890 1570.910 3377.070 ;
        RECT 1569.730 3374.290 1570.910 3375.470 ;
        RECT 1569.730 3195.890 1570.910 3197.070 ;
        RECT 1569.730 3194.290 1570.910 3195.470 ;
        RECT 1569.730 3015.890 1570.910 3017.070 ;
        RECT 1569.730 3014.290 1570.910 3015.470 ;
        RECT 1569.730 2835.890 1570.910 2837.070 ;
        RECT 1569.730 2834.290 1570.910 2835.470 ;
        RECT 1569.730 2655.890 1570.910 2657.070 ;
        RECT 1569.730 2654.290 1570.910 2655.470 ;
        RECT 1569.730 2475.890 1570.910 2477.070 ;
        RECT 1569.730 2474.290 1570.910 2475.470 ;
        RECT 1569.730 2295.890 1570.910 2297.070 ;
        RECT 1569.730 2294.290 1570.910 2295.470 ;
        RECT 1569.730 2115.890 1570.910 2117.070 ;
        RECT 1569.730 2114.290 1570.910 2115.470 ;
        RECT 1569.730 1935.890 1570.910 1937.070 ;
        RECT 1569.730 1934.290 1570.910 1935.470 ;
        RECT 1569.730 1755.890 1570.910 1757.070 ;
        RECT 1569.730 1754.290 1570.910 1755.470 ;
        RECT 1569.730 1575.890 1570.910 1577.070 ;
        RECT 1569.730 1574.290 1570.910 1575.470 ;
        RECT 1569.730 1395.890 1570.910 1397.070 ;
        RECT 1569.730 1394.290 1570.910 1395.470 ;
        RECT 1569.730 1215.890 1570.910 1217.070 ;
        RECT 1569.730 1214.290 1570.910 1215.470 ;
        RECT 1569.730 1035.890 1570.910 1037.070 ;
        RECT 1569.730 1034.290 1570.910 1035.470 ;
        RECT 1569.730 855.890 1570.910 857.070 ;
        RECT 1569.730 854.290 1570.910 855.470 ;
        RECT 1569.730 675.890 1570.910 677.070 ;
        RECT 1569.730 674.290 1570.910 675.470 ;
        RECT 1569.730 495.890 1570.910 497.070 ;
        RECT 1569.730 494.290 1570.910 495.470 ;
        RECT 1569.730 315.890 1570.910 317.070 ;
        RECT 1569.730 314.290 1570.910 315.470 ;
        RECT 1569.730 135.890 1570.910 137.070 ;
        RECT 1569.730 134.290 1570.910 135.470 ;
        RECT 1569.730 -25.910 1570.910 -24.730 ;
        RECT 1569.730 -27.510 1570.910 -26.330 ;
        RECT 1749.730 3546.010 1750.910 3547.190 ;
        RECT 1749.730 3544.410 1750.910 3545.590 ;
        RECT 1749.730 3375.890 1750.910 3377.070 ;
        RECT 1749.730 3374.290 1750.910 3375.470 ;
        RECT 1749.730 3195.890 1750.910 3197.070 ;
        RECT 1749.730 3194.290 1750.910 3195.470 ;
        RECT 1749.730 3015.890 1750.910 3017.070 ;
        RECT 1749.730 3014.290 1750.910 3015.470 ;
        RECT 1749.730 2835.890 1750.910 2837.070 ;
        RECT 1749.730 2834.290 1750.910 2835.470 ;
        RECT 1749.730 2655.890 1750.910 2657.070 ;
        RECT 1749.730 2654.290 1750.910 2655.470 ;
        RECT 1749.730 2475.890 1750.910 2477.070 ;
        RECT 1749.730 2474.290 1750.910 2475.470 ;
        RECT 1749.730 2295.890 1750.910 2297.070 ;
        RECT 1749.730 2294.290 1750.910 2295.470 ;
        RECT 1749.730 2115.890 1750.910 2117.070 ;
        RECT 1749.730 2114.290 1750.910 2115.470 ;
        RECT 1749.730 1935.890 1750.910 1937.070 ;
        RECT 1749.730 1934.290 1750.910 1935.470 ;
        RECT 1749.730 1755.890 1750.910 1757.070 ;
        RECT 1749.730 1754.290 1750.910 1755.470 ;
        RECT 1749.730 1575.890 1750.910 1577.070 ;
        RECT 1749.730 1574.290 1750.910 1575.470 ;
        RECT 1749.730 1395.890 1750.910 1397.070 ;
        RECT 1749.730 1394.290 1750.910 1395.470 ;
        RECT 1749.730 1215.890 1750.910 1217.070 ;
        RECT 1749.730 1214.290 1750.910 1215.470 ;
        RECT 1749.730 1035.890 1750.910 1037.070 ;
        RECT 1749.730 1034.290 1750.910 1035.470 ;
        RECT 1749.730 855.890 1750.910 857.070 ;
        RECT 1749.730 854.290 1750.910 855.470 ;
        RECT 1749.730 675.890 1750.910 677.070 ;
        RECT 1749.730 674.290 1750.910 675.470 ;
        RECT 1749.730 495.890 1750.910 497.070 ;
        RECT 1749.730 494.290 1750.910 495.470 ;
        RECT 1749.730 315.890 1750.910 317.070 ;
        RECT 1749.730 314.290 1750.910 315.470 ;
        RECT 1749.730 135.890 1750.910 137.070 ;
        RECT 1749.730 134.290 1750.910 135.470 ;
        RECT 1749.730 -25.910 1750.910 -24.730 ;
        RECT 1749.730 -27.510 1750.910 -26.330 ;
        RECT 1929.730 3546.010 1930.910 3547.190 ;
        RECT 1929.730 3544.410 1930.910 3545.590 ;
        RECT 1929.730 3375.890 1930.910 3377.070 ;
        RECT 1929.730 3374.290 1930.910 3375.470 ;
        RECT 1929.730 3195.890 1930.910 3197.070 ;
        RECT 1929.730 3194.290 1930.910 3195.470 ;
        RECT 1929.730 3015.890 1930.910 3017.070 ;
        RECT 1929.730 3014.290 1930.910 3015.470 ;
        RECT 1929.730 2835.890 1930.910 2837.070 ;
        RECT 1929.730 2834.290 1930.910 2835.470 ;
        RECT 1929.730 2655.890 1930.910 2657.070 ;
        RECT 1929.730 2654.290 1930.910 2655.470 ;
        RECT 1929.730 2475.890 1930.910 2477.070 ;
        RECT 1929.730 2474.290 1930.910 2475.470 ;
        RECT 1929.730 2295.890 1930.910 2297.070 ;
        RECT 1929.730 2294.290 1930.910 2295.470 ;
        RECT 1929.730 2115.890 1930.910 2117.070 ;
        RECT 1929.730 2114.290 1930.910 2115.470 ;
        RECT 1929.730 1935.890 1930.910 1937.070 ;
        RECT 1929.730 1934.290 1930.910 1935.470 ;
        RECT 1929.730 1755.890 1930.910 1757.070 ;
        RECT 1929.730 1754.290 1930.910 1755.470 ;
        RECT 1929.730 1575.890 1930.910 1577.070 ;
        RECT 1929.730 1574.290 1930.910 1575.470 ;
        RECT 1929.730 1395.890 1930.910 1397.070 ;
        RECT 1929.730 1394.290 1930.910 1395.470 ;
        RECT 1929.730 1215.890 1930.910 1217.070 ;
        RECT 1929.730 1214.290 1930.910 1215.470 ;
        RECT 1929.730 1035.890 1930.910 1037.070 ;
        RECT 1929.730 1034.290 1930.910 1035.470 ;
        RECT 1929.730 855.890 1930.910 857.070 ;
        RECT 1929.730 854.290 1930.910 855.470 ;
        RECT 1929.730 675.890 1930.910 677.070 ;
        RECT 1929.730 674.290 1930.910 675.470 ;
        RECT 1929.730 495.890 1930.910 497.070 ;
        RECT 1929.730 494.290 1930.910 495.470 ;
        RECT 1929.730 315.890 1930.910 317.070 ;
        RECT 1929.730 314.290 1930.910 315.470 ;
        RECT 1929.730 135.890 1930.910 137.070 ;
        RECT 1929.730 134.290 1930.910 135.470 ;
        RECT 1929.730 -25.910 1930.910 -24.730 ;
        RECT 1929.730 -27.510 1930.910 -26.330 ;
        RECT 2109.730 3546.010 2110.910 3547.190 ;
        RECT 2109.730 3544.410 2110.910 3545.590 ;
        RECT 2109.730 3375.890 2110.910 3377.070 ;
        RECT 2109.730 3374.290 2110.910 3375.470 ;
        RECT 2109.730 3195.890 2110.910 3197.070 ;
        RECT 2109.730 3194.290 2110.910 3195.470 ;
        RECT 2109.730 3015.890 2110.910 3017.070 ;
        RECT 2109.730 3014.290 2110.910 3015.470 ;
        RECT 2109.730 2835.890 2110.910 2837.070 ;
        RECT 2109.730 2834.290 2110.910 2835.470 ;
        RECT 2109.730 2655.890 2110.910 2657.070 ;
        RECT 2109.730 2654.290 2110.910 2655.470 ;
        RECT 2109.730 2475.890 2110.910 2477.070 ;
        RECT 2109.730 2474.290 2110.910 2475.470 ;
        RECT 2109.730 2295.890 2110.910 2297.070 ;
        RECT 2109.730 2294.290 2110.910 2295.470 ;
        RECT 2109.730 2115.890 2110.910 2117.070 ;
        RECT 2109.730 2114.290 2110.910 2115.470 ;
        RECT 2109.730 1935.890 2110.910 1937.070 ;
        RECT 2109.730 1934.290 2110.910 1935.470 ;
        RECT 2109.730 1755.890 2110.910 1757.070 ;
        RECT 2109.730 1754.290 2110.910 1755.470 ;
        RECT 2109.730 1575.890 2110.910 1577.070 ;
        RECT 2109.730 1574.290 2110.910 1575.470 ;
        RECT 2109.730 1395.890 2110.910 1397.070 ;
        RECT 2109.730 1394.290 2110.910 1395.470 ;
        RECT 2109.730 1215.890 2110.910 1217.070 ;
        RECT 2109.730 1214.290 2110.910 1215.470 ;
        RECT 2109.730 1035.890 2110.910 1037.070 ;
        RECT 2109.730 1034.290 2110.910 1035.470 ;
        RECT 2109.730 855.890 2110.910 857.070 ;
        RECT 2109.730 854.290 2110.910 855.470 ;
        RECT 2109.730 675.890 2110.910 677.070 ;
        RECT 2109.730 674.290 2110.910 675.470 ;
        RECT 2109.730 495.890 2110.910 497.070 ;
        RECT 2109.730 494.290 2110.910 495.470 ;
        RECT 2109.730 315.890 2110.910 317.070 ;
        RECT 2109.730 314.290 2110.910 315.470 ;
        RECT 2109.730 135.890 2110.910 137.070 ;
        RECT 2109.730 134.290 2110.910 135.470 ;
        RECT 2109.730 -25.910 2110.910 -24.730 ;
        RECT 2109.730 -27.510 2110.910 -26.330 ;
        RECT 2289.730 3546.010 2290.910 3547.190 ;
        RECT 2289.730 3544.410 2290.910 3545.590 ;
        RECT 2289.730 3375.890 2290.910 3377.070 ;
        RECT 2289.730 3374.290 2290.910 3375.470 ;
        RECT 2289.730 3195.890 2290.910 3197.070 ;
        RECT 2289.730 3194.290 2290.910 3195.470 ;
        RECT 2289.730 3015.890 2290.910 3017.070 ;
        RECT 2289.730 3014.290 2290.910 3015.470 ;
        RECT 2289.730 2835.890 2290.910 2837.070 ;
        RECT 2289.730 2834.290 2290.910 2835.470 ;
        RECT 2289.730 2655.890 2290.910 2657.070 ;
        RECT 2289.730 2654.290 2290.910 2655.470 ;
        RECT 2289.730 2475.890 2290.910 2477.070 ;
        RECT 2289.730 2474.290 2290.910 2475.470 ;
        RECT 2289.730 2295.890 2290.910 2297.070 ;
        RECT 2289.730 2294.290 2290.910 2295.470 ;
        RECT 2289.730 2115.890 2290.910 2117.070 ;
        RECT 2289.730 2114.290 2290.910 2115.470 ;
        RECT 2289.730 1935.890 2290.910 1937.070 ;
        RECT 2289.730 1934.290 2290.910 1935.470 ;
        RECT 2289.730 1755.890 2290.910 1757.070 ;
        RECT 2289.730 1754.290 2290.910 1755.470 ;
        RECT 2289.730 1575.890 2290.910 1577.070 ;
        RECT 2289.730 1574.290 2290.910 1575.470 ;
        RECT 2289.730 1395.890 2290.910 1397.070 ;
        RECT 2289.730 1394.290 2290.910 1395.470 ;
        RECT 2289.730 1215.890 2290.910 1217.070 ;
        RECT 2289.730 1214.290 2290.910 1215.470 ;
        RECT 2289.730 1035.890 2290.910 1037.070 ;
        RECT 2289.730 1034.290 2290.910 1035.470 ;
        RECT 2289.730 855.890 2290.910 857.070 ;
        RECT 2289.730 854.290 2290.910 855.470 ;
        RECT 2289.730 675.890 2290.910 677.070 ;
        RECT 2289.730 674.290 2290.910 675.470 ;
        RECT 2289.730 495.890 2290.910 497.070 ;
        RECT 2289.730 494.290 2290.910 495.470 ;
        RECT 2289.730 315.890 2290.910 317.070 ;
        RECT 2289.730 314.290 2290.910 315.470 ;
        RECT 2289.730 135.890 2290.910 137.070 ;
        RECT 2289.730 134.290 2290.910 135.470 ;
        RECT 2289.730 -25.910 2290.910 -24.730 ;
        RECT 2289.730 -27.510 2290.910 -26.330 ;
        RECT 2469.730 3546.010 2470.910 3547.190 ;
        RECT 2469.730 3544.410 2470.910 3545.590 ;
        RECT 2469.730 3375.890 2470.910 3377.070 ;
        RECT 2469.730 3374.290 2470.910 3375.470 ;
        RECT 2469.730 3195.890 2470.910 3197.070 ;
        RECT 2469.730 3194.290 2470.910 3195.470 ;
        RECT 2469.730 3015.890 2470.910 3017.070 ;
        RECT 2469.730 3014.290 2470.910 3015.470 ;
        RECT 2469.730 2835.890 2470.910 2837.070 ;
        RECT 2469.730 2834.290 2470.910 2835.470 ;
        RECT 2469.730 2655.890 2470.910 2657.070 ;
        RECT 2469.730 2654.290 2470.910 2655.470 ;
        RECT 2469.730 2475.890 2470.910 2477.070 ;
        RECT 2469.730 2474.290 2470.910 2475.470 ;
        RECT 2469.730 2295.890 2470.910 2297.070 ;
        RECT 2469.730 2294.290 2470.910 2295.470 ;
        RECT 2469.730 2115.890 2470.910 2117.070 ;
        RECT 2469.730 2114.290 2470.910 2115.470 ;
        RECT 2469.730 1935.890 2470.910 1937.070 ;
        RECT 2469.730 1934.290 2470.910 1935.470 ;
        RECT 2469.730 1755.890 2470.910 1757.070 ;
        RECT 2469.730 1754.290 2470.910 1755.470 ;
        RECT 2469.730 1575.890 2470.910 1577.070 ;
        RECT 2469.730 1574.290 2470.910 1575.470 ;
        RECT 2469.730 1395.890 2470.910 1397.070 ;
        RECT 2469.730 1394.290 2470.910 1395.470 ;
        RECT 2469.730 1215.890 2470.910 1217.070 ;
        RECT 2469.730 1214.290 2470.910 1215.470 ;
        RECT 2469.730 1035.890 2470.910 1037.070 ;
        RECT 2469.730 1034.290 2470.910 1035.470 ;
        RECT 2469.730 855.890 2470.910 857.070 ;
        RECT 2469.730 854.290 2470.910 855.470 ;
        RECT 2469.730 675.890 2470.910 677.070 ;
        RECT 2469.730 674.290 2470.910 675.470 ;
        RECT 2469.730 495.890 2470.910 497.070 ;
        RECT 2469.730 494.290 2470.910 495.470 ;
        RECT 2469.730 315.890 2470.910 317.070 ;
        RECT 2469.730 314.290 2470.910 315.470 ;
        RECT 2469.730 135.890 2470.910 137.070 ;
        RECT 2469.730 134.290 2470.910 135.470 ;
        RECT 2469.730 -25.910 2470.910 -24.730 ;
        RECT 2469.730 -27.510 2470.910 -26.330 ;
        RECT 2649.730 3546.010 2650.910 3547.190 ;
        RECT 2649.730 3544.410 2650.910 3545.590 ;
        RECT 2649.730 3375.890 2650.910 3377.070 ;
        RECT 2649.730 3374.290 2650.910 3375.470 ;
        RECT 2649.730 3195.890 2650.910 3197.070 ;
        RECT 2649.730 3194.290 2650.910 3195.470 ;
        RECT 2649.730 3015.890 2650.910 3017.070 ;
        RECT 2649.730 3014.290 2650.910 3015.470 ;
        RECT 2649.730 2835.890 2650.910 2837.070 ;
        RECT 2649.730 2834.290 2650.910 2835.470 ;
        RECT 2649.730 2655.890 2650.910 2657.070 ;
        RECT 2649.730 2654.290 2650.910 2655.470 ;
        RECT 2649.730 2475.890 2650.910 2477.070 ;
        RECT 2649.730 2474.290 2650.910 2475.470 ;
        RECT 2649.730 2295.890 2650.910 2297.070 ;
        RECT 2649.730 2294.290 2650.910 2295.470 ;
        RECT 2649.730 2115.890 2650.910 2117.070 ;
        RECT 2649.730 2114.290 2650.910 2115.470 ;
        RECT 2649.730 1935.890 2650.910 1937.070 ;
        RECT 2649.730 1934.290 2650.910 1935.470 ;
        RECT 2649.730 1755.890 2650.910 1757.070 ;
        RECT 2649.730 1754.290 2650.910 1755.470 ;
        RECT 2649.730 1575.890 2650.910 1577.070 ;
        RECT 2649.730 1574.290 2650.910 1575.470 ;
        RECT 2649.730 1395.890 2650.910 1397.070 ;
        RECT 2649.730 1394.290 2650.910 1395.470 ;
        RECT 2649.730 1215.890 2650.910 1217.070 ;
        RECT 2649.730 1214.290 2650.910 1215.470 ;
        RECT 2649.730 1035.890 2650.910 1037.070 ;
        RECT 2649.730 1034.290 2650.910 1035.470 ;
        RECT 2649.730 855.890 2650.910 857.070 ;
        RECT 2649.730 854.290 2650.910 855.470 ;
        RECT 2649.730 675.890 2650.910 677.070 ;
        RECT 2649.730 674.290 2650.910 675.470 ;
        RECT 2649.730 495.890 2650.910 497.070 ;
        RECT 2649.730 494.290 2650.910 495.470 ;
        RECT 2649.730 315.890 2650.910 317.070 ;
        RECT 2649.730 314.290 2650.910 315.470 ;
        RECT 2649.730 135.890 2650.910 137.070 ;
        RECT 2649.730 134.290 2650.910 135.470 ;
        RECT 2649.730 -25.910 2650.910 -24.730 ;
        RECT 2649.730 -27.510 2650.910 -26.330 ;
        RECT 2829.730 3546.010 2830.910 3547.190 ;
        RECT 2829.730 3544.410 2830.910 3545.590 ;
        RECT 2829.730 3375.890 2830.910 3377.070 ;
        RECT 2829.730 3374.290 2830.910 3375.470 ;
        RECT 2829.730 3195.890 2830.910 3197.070 ;
        RECT 2829.730 3194.290 2830.910 3195.470 ;
        RECT 2829.730 3015.890 2830.910 3017.070 ;
        RECT 2829.730 3014.290 2830.910 3015.470 ;
        RECT 2829.730 2835.890 2830.910 2837.070 ;
        RECT 2829.730 2834.290 2830.910 2835.470 ;
        RECT 2829.730 2655.890 2830.910 2657.070 ;
        RECT 2829.730 2654.290 2830.910 2655.470 ;
        RECT 2829.730 2475.890 2830.910 2477.070 ;
        RECT 2829.730 2474.290 2830.910 2475.470 ;
        RECT 2829.730 2295.890 2830.910 2297.070 ;
        RECT 2829.730 2294.290 2830.910 2295.470 ;
        RECT 2829.730 2115.890 2830.910 2117.070 ;
        RECT 2829.730 2114.290 2830.910 2115.470 ;
        RECT 2829.730 1935.890 2830.910 1937.070 ;
        RECT 2829.730 1934.290 2830.910 1935.470 ;
        RECT 2829.730 1755.890 2830.910 1757.070 ;
        RECT 2829.730 1754.290 2830.910 1755.470 ;
        RECT 2829.730 1575.890 2830.910 1577.070 ;
        RECT 2829.730 1574.290 2830.910 1575.470 ;
        RECT 2829.730 1395.890 2830.910 1397.070 ;
        RECT 2829.730 1394.290 2830.910 1395.470 ;
        RECT 2829.730 1215.890 2830.910 1217.070 ;
        RECT 2829.730 1214.290 2830.910 1215.470 ;
        RECT 2829.730 1035.890 2830.910 1037.070 ;
        RECT 2829.730 1034.290 2830.910 1035.470 ;
        RECT 2829.730 855.890 2830.910 857.070 ;
        RECT 2829.730 854.290 2830.910 855.470 ;
        RECT 2829.730 675.890 2830.910 677.070 ;
        RECT 2829.730 674.290 2830.910 675.470 ;
        RECT 2829.730 495.890 2830.910 497.070 ;
        RECT 2829.730 494.290 2830.910 495.470 ;
        RECT 2829.730 315.890 2830.910 317.070 ;
        RECT 2829.730 314.290 2830.910 315.470 ;
        RECT 2829.730 135.890 2830.910 137.070 ;
        RECT 2829.730 134.290 2830.910 135.470 ;
        RECT 2829.730 -25.910 2830.910 -24.730 ;
        RECT 2829.730 -27.510 2830.910 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3375.890 2951.690 3377.070 ;
        RECT 2950.510 3374.290 2951.690 3375.470 ;
        RECT 2950.510 3195.890 2951.690 3197.070 ;
        RECT 2950.510 3194.290 2951.690 3195.470 ;
        RECT 2950.510 3015.890 2951.690 3017.070 ;
        RECT 2950.510 3014.290 2951.690 3015.470 ;
        RECT 2950.510 2835.890 2951.690 2837.070 ;
        RECT 2950.510 2834.290 2951.690 2835.470 ;
        RECT 2950.510 2655.890 2951.690 2657.070 ;
        RECT 2950.510 2654.290 2951.690 2655.470 ;
        RECT 2950.510 2475.890 2951.690 2477.070 ;
        RECT 2950.510 2474.290 2951.690 2475.470 ;
        RECT 2950.510 2295.890 2951.690 2297.070 ;
        RECT 2950.510 2294.290 2951.690 2295.470 ;
        RECT 2950.510 2115.890 2951.690 2117.070 ;
        RECT 2950.510 2114.290 2951.690 2115.470 ;
        RECT 2950.510 1935.890 2951.690 1937.070 ;
        RECT 2950.510 1934.290 2951.690 1935.470 ;
        RECT 2950.510 1755.890 2951.690 1757.070 ;
        RECT 2950.510 1754.290 2951.690 1755.470 ;
        RECT 2950.510 1575.890 2951.690 1577.070 ;
        RECT 2950.510 1574.290 2951.690 1575.470 ;
        RECT 2950.510 1395.890 2951.690 1397.070 ;
        RECT 2950.510 1394.290 2951.690 1395.470 ;
        RECT 2950.510 1215.890 2951.690 1217.070 ;
        RECT 2950.510 1214.290 2951.690 1215.470 ;
        RECT 2950.510 1035.890 2951.690 1037.070 ;
        RECT 2950.510 1034.290 2951.690 1035.470 ;
        RECT 2950.510 855.890 2951.690 857.070 ;
        RECT 2950.510 854.290 2951.690 855.470 ;
        RECT 2950.510 675.890 2951.690 677.070 ;
        RECT 2950.510 674.290 2951.690 675.470 ;
        RECT 2950.510 495.890 2951.690 497.070 ;
        RECT 2950.510 494.290 2951.690 495.470 ;
        RECT 2950.510 315.890 2951.690 317.070 ;
        RECT 2950.510 314.290 2951.690 315.470 ;
        RECT 2950.510 135.890 2951.690 137.070 ;
        RECT 2950.510 134.290 2951.690 135.470 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.930 3547.250 -30.030 3547.310 ;
        RECT 128.870 3547.250 131.770 3547.310 ;
        RECT 308.870 3547.250 311.770 3547.310 ;
        RECT 488.870 3547.250 491.770 3547.310 ;
        RECT 668.870 3547.250 671.770 3547.310 ;
        RECT 848.870 3547.250 851.770 3547.310 ;
        RECT 1028.870 3547.250 1031.770 3547.310 ;
        RECT 1208.870 3547.250 1211.770 3547.310 ;
        RECT 1388.870 3547.250 1391.770 3547.310 ;
        RECT 1568.870 3547.250 1571.770 3547.310 ;
        RECT 1748.870 3547.250 1751.770 3547.310 ;
        RECT 1928.870 3547.250 1931.770 3547.310 ;
        RECT 2108.870 3547.250 2111.770 3547.310 ;
        RECT 2288.870 3547.250 2291.770 3547.310 ;
        RECT 2468.870 3547.250 2471.770 3547.310 ;
        RECT 2648.870 3547.250 2651.770 3547.310 ;
        RECT 2828.870 3547.250 2831.770 3547.310 ;
        RECT 2949.650 3547.250 2952.550 3547.310 ;
        RECT -32.930 3544.350 2952.550 3547.250 ;
        RECT -32.930 3544.290 -30.030 3544.350 ;
        RECT 128.870 3544.290 131.770 3544.350 ;
        RECT 308.870 3544.290 311.770 3544.350 ;
        RECT 488.870 3544.290 491.770 3544.350 ;
        RECT 668.870 3544.290 671.770 3544.350 ;
        RECT 848.870 3544.290 851.770 3544.350 ;
        RECT 1028.870 3544.290 1031.770 3544.350 ;
        RECT 1208.870 3544.290 1211.770 3544.350 ;
        RECT 1388.870 3544.290 1391.770 3544.350 ;
        RECT 1568.870 3544.290 1571.770 3544.350 ;
        RECT 1748.870 3544.290 1751.770 3544.350 ;
        RECT 1928.870 3544.290 1931.770 3544.350 ;
        RECT 2108.870 3544.290 2111.770 3544.350 ;
        RECT 2288.870 3544.290 2291.770 3544.350 ;
        RECT 2468.870 3544.290 2471.770 3544.350 ;
        RECT 2648.870 3544.290 2651.770 3544.350 ;
        RECT 2828.870 3544.290 2831.770 3544.350 ;
        RECT 2949.650 3544.290 2952.550 3544.350 ;
        RECT -32.930 3377.130 -30.030 3377.190 ;
        RECT 128.870 3377.130 131.770 3377.190 ;
        RECT 308.870 3377.130 311.770 3377.190 ;
        RECT 488.870 3377.130 491.770 3377.190 ;
        RECT 668.870 3377.130 671.770 3377.190 ;
        RECT 848.870 3377.130 851.770 3377.190 ;
        RECT 1028.870 3377.130 1031.770 3377.190 ;
        RECT 1208.870 3377.130 1211.770 3377.190 ;
        RECT 1388.870 3377.130 1391.770 3377.190 ;
        RECT 1568.870 3377.130 1571.770 3377.190 ;
        RECT 1748.870 3377.130 1751.770 3377.190 ;
        RECT 1928.870 3377.130 1931.770 3377.190 ;
        RECT 2108.870 3377.130 2111.770 3377.190 ;
        RECT 2288.870 3377.130 2291.770 3377.190 ;
        RECT 2468.870 3377.130 2471.770 3377.190 ;
        RECT 2648.870 3377.130 2651.770 3377.190 ;
        RECT 2828.870 3377.130 2831.770 3377.190 ;
        RECT 2949.650 3377.130 2952.550 3377.190 ;
        RECT -32.930 3374.230 2952.550 3377.130 ;
        RECT -32.930 3374.170 -30.030 3374.230 ;
        RECT 128.870 3374.170 131.770 3374.230 ;
        RECT 308.870 3374.170 311.770 3374.230 ;
        RECT 488.870 3374.170 491.770 3374.230 ;
        RECT 668.870 3374.170 671.770 3374.230 ;
        RECT 848.870 3374.170 851.770 3374.230 ;
        RECT 1028.870 3374.170 1031.770 3374.230 ;
        RECT 1208.870 3374.170 1211.770 3374.230 ;
        RECT 1388.870 3374.170 1391.770 3374.230 ;
        RECT 1568.870 3374.170 1571.770 3374.230 ;
        RECT 1748.870 3374.170 1751.770 3374.230 ;
        RECT 1928.870 3374.170 1931.770 3374.230 ;
        RECT 2108.870 3374.170 2111.770 3374.230 ;
        RECT 2288.870 3374.170 2291.770 3374.230 ;
        RECT 2468.870 3374.170 2471.770 3374.230 ;
        RECT 2648.870 3374.170 2651.770 3374.230 ;
        RECT 2828.870 3374.170 2831.770 3374.230 ;
        RECT 2949.650 3374.170 2952.550 3374.230 ;
        RECT -32.930 3197.130 -30.030 3197.190 ;
        RECT 128.870 3197.130 131.770 3197.190 ;
        RECT 308.870 3197.130 311.770 3197.190 ;
        RECT 488.870 3197.130 491.770 3197.190 ;
        RECT 668.870 3197.130 671.770 3197.190 ;
        RECT 848.870 3197.130 851.770 3197.190 ;
        RECT 1028.870 3197.130 1031.770 3197.190 ;
        RECT 1208.870 3197.130 1211.770 3197.190 ;
        RECT 1388.870 3197.130 1391.770 3197.190 ;
        RECT 1568.870 3197.130 1571.770 3197.190 ;
        RECT 1748.870 3197.130 1751.770 3197.190 ;
        RECT 1928.870 3197.130 1931.770 3197.190 ;
        RECT 2108.870 3197.130 2111.770 3197.190 ;
        RECT 2288.870 3197.130 2291.770 3197.190 ;
        RECT 2468.870 3197.130 2471.770 3197.190 ;
        RECT 2648.870 3197.130 2651.770 3197.190 ;
        RECT 2828.870 3197.130 2831.770 3197.190 ;
        RECT 2949.650 3197.130 2952.550 3197.190 ;
        RECT -32.930 3194.230 2952.550 3197.130 ;
        RECT -32.930 3194.170 -30.030 3194.230 ;
        RECT 128.870 3194.170 131.770 3194.230 ;
        RECT 308.870 3194.170 311.770 3194.230 ;
        RECT 488.870 3194.170 491.770 3194.230 ;
        RECT 668.870 3194.170 671.770 3194.230 ;
        RECT 848.870 3194.170 851.770 3194.230 ;
        RECT 1028.870 3194.170 1031.770 3194.230 ;
        RECT 1208.870 3194.170 1211.770 3194.230 ;
        RECT 1388.870 3194.170 1391.770 3194.230 ;
        RECT 1568.870 3194.170 1571.770 3194.230 ;
        RECT 1748.870 3194.170 1751.770 3194.230 ;
        RECT 1928.870 3194.170 1931.770 3194.230 ;
        RECT 2108.870 3194.170 2111.770 3194.230 ;
        RECT 2288.870 3194.170 2291.770 3194.230 ;
        RECT 2468.870 3194.170 2471.770 3194.230 ;
        RECT 2648.870 3194.170 2651.770 3194.230 ;
        RECT 2828.870 3194.170 2831.770 3194.230 ;
        RECT 2949.650 3194.170 2952.550 3194.230 ;
        RECT -32.930 3017.130 -30.030 3017.190 ;
        RECT 128.870 3017.130 131.770 3017.190 ;
        RECT 308.870 3017.130 311.770 3017.190 ;
        RECT 488.870 3017.130 491.770 3017.190 ;
        RECT 668.870 3017.130 671.770 3017.190 ;
        RECT 848.870 3017.130 851.770 3017.190 ;
        RECT 1028.870 3017.130 1031.770 3017.190 ;
        RECT 1208.870 3017.130 1211.770 3017.190 ;
        RECT 1388.870 3017.130 1391.770 3017.190 ;
        RECT 1568.870 3017.130 1571.770 3017.190 ;
        RECT 1748.870 3017.130 1751.770 3017.190 ;
        RECT 1928.870 3017.130 1931.770 3017.190 ;
        RECT 2108.870 3017.130 2111.770 3017.190 ;
        RECT 2288.870 3017.130 2291.770 3017.190 ;
        RECT 2468.870 3017.130 2471.770 3017.190 ;
        RECT 2648.870 3017.130 2651.770 3017.190 ;
        RECT 2828.870 3017.130 2831.770 3017.190 ;
        RECT 2949.650 3017.130 2952.550 3017.190 ;
        RECT -32.930 3014.230 2952.550 3017.130 ;
        RECT -32.930 3014.170 -30.030 3014.230 ;
        RECT 128.870 3014.170 131.770 3014.230 ;
        RECT 308.870 3014.170 311.770 3014.230 ;
        RECT 488.870 3014.170 491.770 3014.230 ;
        RECT 668.870 3014.170 671.770 3014.230 ;
        RECT 848.870 3014.170 851.770 3014.230 ;
        RECT 1028.870 3014.170 1031.770 3014.230 ;
        RECT 1208.870 3014.170 1211.770 3014.230 ;
        RECT 1388.870 3014.170 1391.770 3014.230 ;
        RECT 1568.870 3014.170 1571.770 3014.230 ;
        RECT 1748.870 3014.170 1751.770 3014.230 ;
        RECT 1928.870 3014.170 1931.770 3014.230 ;
        RECT 2108.870 3014.170 2111.770 3014.230 ;
        RECT 2288.870 3014.170 2291.770 3014.230 ;
        RECT 2468.870 3014.170 2471.770 3014.230 ;
        RECT 2648.870 3014.170 2651.770 3014.230 ;
        RECT 2828.870 3014.170 2831.770 3014.230 ;
        RECT 2949.650 3014.170 2952.550 3014.230 ;
        RECT -32.930 2837.130 -30.030 2837.190 ;
        RECT 128.870 2837.130 131.770 2837.190 ;
        RECT 308.870 2837.130 311.770 2837.190 ;
        RECT 488.870 2837.130 491.770 2837.190 ;
        RECT 668.870 2837.130 671.770 2837.190 ;
        RECT 848.870 2837.130 851.770 2837.190 ;
        RECT 1028.870 2837.130 1031.770 2837.190 ;
        RECT 1208.870 2837.130 1211.770 2837.190 ;
        RECT 1388.870 2837.130 1391.770 2837.190 ;
        RECT 1568.870 2837.130 1571.770 2837.190 ;
        RECT 1748.870 2837.130 1751.770 2837.190 ;
        RECT 1928.870 2837.130 1931.770 2837.190 ;
        RECT 2108.870 2837.130 2111.770 2837.190 ;
        RECT 2288.870 2837.130 2291.770 2837.190 ;
        RECT 2468.870 2837.130 2471.770 2837.190 ;
        RECT 2648.870 2837.130 2651.770 2837.190 ;
        RECT 2828.870 2837.130 2831.770 2837.190 ;
        RECT 2949.650 2837.130 2952.550 2837.190 ;
        RECT -32.930 2834.230 2952.550 2837.130 ;
        RECT -32.930 2834.170 -30.030 2834.230 ;
        RECT 128.870 2834.170 131.770 2834.230 ;
        RECT 308.870 2834.170 311.770 2834.230 ;
        RECT 488.870 2834.170 491.770 2834.230 ;
        RECT 668.870 2834.170 671.770 2834.230 ;
        RECT 848.870 2834.170 851.770 2834.230 ;
        RECT 1028.870 2834.170 1031.770 2834.230 ;
        RECT 1208.870 2834.170 1211.770 2834.230 ;
        RECT 1388.870 2834.170 1391.770 2834.230 ;
        RECT 1568.870 2834.170 1571.770 2834.230 ;
        RECT 1748.870 2834.170 1751.770 2834.230 ;
        RECT 1928.870 2834.170 1931.770 2834.230 ;
        RECT 2108.870 2834.170 2111.770 2834.230 ;
        RECT 2288.870 2834.170 2291.770 2834.230 ;
        RECT 2468.870 2834.170 2471.770 2834.230 ;
        RECT 2648.870 2834.170 2651.770 2834.230 ;
        RECT 2828.870 2834.170 2831.770 2834.230 ;
        RECT 2949.650 2834.170 2952.550 2834.230 ;
        RECT -32.930 2657.130 -30.030 2657.190 ;
        RECT 128.870 2657.130 131.770 2657.190 ;
        RECT 308.870 2657.130 311.770 2657.190 ;
        RECT 488.870 2657.130 491.770 2657.190 ;
        RECT 668.870 2657.130 671.770 2657.190 ;
        RECT 848.870 2657.130 851.770 2657.190 ;
        RECT 1028.870 2657.130 1031.770 2657.190 ;
        RECT 1208.870 2657.130 1211.770 2657.190 ;
        RECT 1388.870 2657.130 1391.770 2657.190 ;
        RECT 1568.870 2657.130 1571.770 2657.190 ;
        RECT 1748.870 2657.130 1751.770 2657.190 ;
        RECT 1928.870 2657.130 1931.770 2657.190 ;
        RECT 2108.870 2657.130 2111.770 2657.190 ;
        RECT 2288.870 2657.130 2291.770 2657.190 ;
        RECT 2468.870 2657.130 2471.770 2657.190 ;
        RECT 2648.870 2657.130 2651.770 2657.190 ;
        RECT 2828.870 2657.130 2831.770 2657.190 ;
        RECT 2949.650 2657.130 2952.550 2657.190 ;
        RECT -32.930 2654.230 2952.550 2657.130 ;
        RECT -32.930 2654.170 -30.030 2654.230 ;
        RECT 128.870 2654.170 131.770 2654.230 ;
        RECT 308.870 2654.170 311.770 2654.230 ;
        RECT 488.870 2654.170 491.770 2654.230 ;
        RECT 668.870 2654.170 671.770 2654.230 ;
        RECT 848.870 2654.170 851.770 2654.230 ;
        RECT 1028.870 2654.170 1031.770 2654.230 ;
        RECT 1208.870 2654.170 1211.770 2654.230 ;
        RECT 1388.870 2654.170 1391.770 2654.230 ;
        RECT 1568.870 2654.170 1571.770 2654.230 ;
        RECT 1748.870 2654.170 1751.770 2654.230 ;
        RECT 1928.870 2654.170 1931.770 2654.230 ;
        RECT 2108.870 2654.170 2111.770 2654.230 ;
        RECT 2288.870 2654.170 2291.770 2654.230 ;
        RECT 2468.870 2654.170 2471.770 2654.230 ;
        RECT 2648.870 2654.170 2651.770 2654.230 ;
        RECT 2828.870 2654.170 2831.770 2654.230 ;
        RECT 2949.650 2654.170 2952.550 2654.230 ;
        RECT -32.930 2477.130 -30.030 2477.190 ;
        RECT 128.870 2477.130 131.770 2477.190 ;
        RECT 308.870 2477.130 311.770 2477.190 ;
        RECT 488.870 2477.130 491.770 2477.190 ;
        RECT 668.870 2477.130 671.770 2477.190 ;
        RECT 848.870 2477.130 851.770 2477.190 ;
        RECT 1028.870 2477.130 1031.770 2477.190 ;
        RECT 1208.870 2477.130 1211.770 2477.190 ;
        RECT 1388.870 2477.130 1391.770 2477.190 ;
        RECT 1568.870 2477.130 1571.770 2477.190 ;
        RECT 1748.870 2477.130 1751.770 2477.190 ;
        RECT 1928.870 2477.130 1931.770 2477.190 ;
        RECT 2108.870 2477.130 2111.770 2477.190 ;
        RECT 2288.870 2477.130 2291.770 2477.190 ;
        RECT 2468.870 2477.130 2471.770 2477.190 ;
        RECT 2648.870 2477.130 2651.770 2477.190 ;
        RECT 2828.870 2477.130 2831.770 2477.190 ;
        RECT 2949.650 2477.130 2952.550 2477.190 ;
        RECT -32.930 2474.230 2952.550 2477.130 ;
        RECT -32.930 2474.170 -30.030 2474.230 ;
        RECT 128.870 2474.170 131.770 2474.230 ;
        RECT 308.870 2474.170 311.770 2474.230 ;
        RECT 488.870 2474.170 491.770 2474.230 ;
        RECT 668.870 2474.170 671.770 2474.230 ;
        RECT 848.870 2474.170 851.770 2474.230 ;
        RECT 1028.870 2474.170 1031.770 2474.230 ;
        RECT 1208.870 2474.170 1211.770 2474.230 ;
        RECT 1388.870 2474.170 1391.770 2474.230 ;
        RECT 1568.870 2474.170 1571.770 2474.230 ;
        RECT 1748.870 2474.170 1751.770 2474.230 ;
        RECT 1928.870 2474.170 1931.770 2474.230 ;
        RECT 2108.870 2474.170 2111.770 2474.230 ;
        RECT 2288.870 2474.170 2291.770 2474.230 ;
        RECT 2468.870 2474.170 2471.770 2474.230 ;
        RECT 2648.870 2474.170 2651.770 2474.230 ;
        RECT 2828.870 2474.170 2831.770 2474.230 ;
        RECT 2949.650 2474.170 2952.550 2474.230 ;
        RECT -32.930 2297.130 -30.030 2297.190 ;
        RECT 128.870 2297.130 131.770 2297.190 ;
        RECT 308.870 2297.130 311.770 2297.190 ;
        RECT 488.870 2297.130 491.770 2297.190 ;
        RECT 668.870 2297.130 671.770 2297.190 ;
        RECT 848.870 2297.130 851.770 2297.190 ;
        RECT 1028.870 2297.130 1031.770 2297.190 ;
        RECT 1208.870 2297.130 1211.770 2297.190 ;
        RECT 1388.870 2297.130 1391.770 2297.190 ;
        RECT 1568.870 2297.130 1571.770 2297.190 ;
        RECT 1748.870 2297.130 1751.770 2297.190 ;
        RECT 1928.870 2297.130 1931.770 2297.190 ;
        RECT 2108.870 2297.130 2111.770 2297.190 ;
        RECT 2288.870 2297.130 2291.770 2297.190 ;
        RECT 2468.870 2297.130 2471.770 2297.190 ;
        RECT 2648.870 2297.130 2651.770 2297.190 ;
        RECT 2828.870 2297.130 2831.770 2297.190 ;
        RECT 2949.650 2297.130 2952.550 2297.190 ;
        RECT -32.930 2294.230 2952.550 2297.130 ;
        RECT -32.930 2294.170 -30.030 2294.230 ;
        RECT 128.870 2294.170 131.770 2294.230 ;
        RECT 308.870 2294.170 311.770 2294.230 ;
        RECT 488.870 2294.170 491.770 2294.230 ;
        RECT 668.870 2294.170 671.770 2294.230 ;
        RECT 848.870 2294.170 851.770 2294.230 ;
        RECT 1028.870 2294.170 1031.770 2294.230 ;
        RECT 1208.870 2294.170 1211.770 2294.230 ;
        RECT 1388.870 2294.170 1391.770 2294.230 ;
        RECT 1568.870 2294.170 1571.770 2294.230 ;
        RECT 1748.870 2294.170 1751.770 2294.230 ;
        RECT 1928.870 2294.170 1931.770 2294.230 ;
        RECT 2108.870 2294.170 2111.770 2294.230 ;
        RECT 2288.870 2294.170 2291.770 2294.230 ;
        RECT 2468.870 2294.170 2471.770 2294.230 ;
        RECT 2648.870 2294.170 2651.770 2294.230 ;
        RECT 2828.870 2294.170 2831.770 2294.230 ;
        RECT 2949.650 2294.170 2952.550 2294.230 ;
        RECT -32.930 2117.130 -30.030 2117.190 ;
        RECT 128.870 2117.130 131.770 2117.190 ;
        RECT 308.870 2117.130 311.770 2117.190 ;
        RECT 488.870 2117.130 491.770 2117.190 ;
        RECT 668.870 2117.130 671.770 2117.190 ;
        RECT 848.870 2117.130 851.770 2117.190 ;
        RECT 1028.870 2117.130 1031.770 2117.190 ;
        RECT 1208.870 2117.130 1211.770 2117.190 ;
        RECT 1388.870 2117.130 1391.770 2117.190 ;
        RECT 1568.870 2117.130 1571.770 2117.190 ;
        RECT 1748.870 2117.130 1751.770 2117.190 ;
        RECT 1928.870 2117.130 1931.770 2117.190 ;
        RECT 2108.870 2117.130 2111.770 2117.190 ;
        RECT 2288.870 2117.130 2291.770 2117.190 ;
        RECT 2468.870 2117.130 2471.770 2117.190 ;
        RECT 2648.870 2117.130 2651.770 2117.190 ;
        RECT 2828.870 2117.130 2831.770 2117.190 ;
        RECT 2949.650 2117.130 2952.550 2117.190 ;
        RECT -32.930 2114.230 2952.550 2117.130 ;
        RECT -32.930 2114.170 -30.030 2114.230 ;
        RECT 128.870 2114.170 131.770 2114.230 ;
        RECT 308.870 2114.170 311.770 2114.230 ;
        RECT 488.870 2114.170 491.770 2114.230 ;
        RECT 668.870 2114.170 671.770 2114.230 ;
        RECT 848.870 2114.170 851.770 2114.230 ;
        RECT 1028.870 2114.170 1031.770 2114.230 ;
        RECT 1208.870 2114.170 1211.770 2114.230 ;
        RECT 1388.870 2114.170 1391.770 2114.230 ;
        RECT 1568.870 2114.170 1571.770 2114.230 ;
        RECT 1748.870 2114.170 1751.770 2114.230 ;
        RECT 1928.870 2114.170 1931.770 2114.230 ;
        RECT 2108.870 2114.170 2111.770 2114.230 ;
        RECT 2288.870 2114.170 2291.770 2114.230 ;
        RECT 2468.870 2114.170 2471.770 2114.230 ;
        RECT 2648.870 2114.170 2651.770 2114.230 ;
        RECT 2828.870 2114.170 2831.770 2114.230 ;
        RECT 2949.650 2114.170 2952.550 2114.230 ;
        RECT -32.930 1937.130 -30.030 1937.190 ;
        RECT 128.870 1937.130 131.770 1937.190 ;
        RECT 308.870 1937.130 311.770 1937.190 ;
        RECT 488.870 1937.130 491.770 1937.190 ;
        RECT 668.870 1937.130 671.770 1937.190 ;
        RECT 848.870 1937.130 851.770 1937.190 ;
        RECT 1028.870 1937.130 1031.770 1937.190 ;
        RECT 1208.870 1937.130 1211.770 1937.190 ;
        RECT 1388.870 1937.130 1391.770 1937.190 ;
        RECT 1568.870 1937.130 1571.770 1937.190 ;
        RECT 1748.870 1937.130 1751.770 1937.190 ;
        RECT 1928.870 1937.130 1931.770 1937.190 ;
        RECT 2108.870 1937.130 2111.770 1937.190 ;
        RECT 2288.870 1937.130 2291.770 1937.190 ;
        RECT 2468.870 1937.130 2471.770 1937.190 ;
        RECT 2648.870 1937.130 2651.770 1937.190 ;
        RECT 2828.870 1937.130 2831.770 1937.190 ;
        RECT 2949.650 1937.130 2952.550 1937.190 ;
        RECT -32.930 1934.230 2952.550 1937.130 ;
        RECT -32.930 1934.170 -30.030 1934.230 ;
        RECT 128.870 1934.170 131.770 1934.230 ;
        RECT 308.870 1934.170 311.770 1934.230 ;
        RECT 488.870 1934.170 491.770 1934.230 ;
        RECT 668.870 1934.170 671.770 1934.230 ;
        RECT 848.870 1934.170 851.770 1934.230 ;
        RECT 1028.870 1934.170 1031.770 1934.230 ;
        RECT 1208.870 1934.170 1211.770 1934.230 ;
        RECT 1388.870 1934.170 1391.770 1934.230 ;
        RECT 1568.870 1934.170 1571.770 1934.230 ;
        RECT 1748.870 1934.170 1751.770 1934.230 ;
        RECT 1928.870 1934.170 1931.770 1934.230 ;
        RECT 2108.870 1934.170 2111.770 1934.230 ;
        RECT 2288.870 1934.170 2291.770 1934.230 ;
        RECT 2468.870 1934.170 2471.770 1934.230 ;
        RECT 2648.870 1934.170 2651.770 1934.230 ;
        RECT 2828.870 1934.170 2831.770 1934.230 ;
        RECT 2949.650 1934.170 2952.550 1934.230 ;
        RECT -32.930 1757.130 -30.030 1757.190 ;
        RECT 128.870 1757.130 131.770 1757.190 ;
        RECT 308.870 1757.130 311.770 1757.190 ;
        RECT 488.870 1757.130 491.770 1757.190 ;
        RECT 668.870 1757.130 671.770 1757.190 ;
        RECT 848.870 1757.130 851.770 1757.190 ;
        RECT 1028.870 1757.130 1031.770 1757.190 ;
        RECT 1208.870 1757.130 1211.770 1757.190 ;
        RECT 1388.870 1757.130 1391.770 1757.190 ;
        RECT 1568.870 1757.130 1571.770 1757.190 ;
        RECT 1748.870 1757.130 1751.770 1757.190 ;
        RECT 1928.870 1757.130 1931.770 1757.190 ;
        RECT 2108.870 1757.130 2111.770 1757.190 ;
        RECT 2288.870 1757.130 2291.770 1757.190 ;
        RECT 2468.870 1757.130 2471.770 1757.190 ;
        RECT 2648.870 1757.130 2651.770 1757.190 ;
        RECT 2828.870 1757.130 2831.770 1757.190 ;
        RECT 2949.650 1757.130 2952.550 1757.190 ;
        RECT -32.930 1754.230 2952.550 1757.130 ;
        RECT -32.930 1754.170 -30.030 1754.230 ;
        RECT 128.870 1754.170 131.770 1754.230 ;
        RECT 308.870 1754.170 311.770 1754.230 ;
        RECT 488.870 1754.170 491.770 1754.230 ;
        RECT 668.870 1754.170 671.770 1754.230 ;
        RECT 848.870 1754.170 851.770 1754.230 ;
        RECT 1028.870 1754.170 1031.770 1754.230 ;
        RECT 1208.870 1754.170 1211.770 1754.230 ;
        RECT 1388.870 1754.170 1391.770 1754.230 ;
        RECT 1568.870 1754.170 1571.770 1754.230 ;
        RECT 1748.870 1754.170 1751.770 1754.230 ;
        RECT 1928.870 1754.170 1931.770 1754.230 ;
        RECT 2108.870 1754.170 2111.770 1754.230 ;
        RECT 2288.870 1754.170 2291.770 1754.230 ;
        RECT 2468.870 1754.170 2471.770 1754.230 ;
        RECT 2648.870 1754.170 2651.770 1754.230 ;
        RECT 2828.870 1754.170 2831.770 1754.230 ;
        RECT 2949.650 1754.170 2952.550 1754.230 ;
        RECT -32.930 1577.130 -30.030 1577.190 ;
        RECT 128.870 1577.130 131.770 1577.190 ;
        RECT 308.870 1577.130 311.770 1577.190 ;
        RECT 488.870 1577.130 491.770 1577.190 ;
        RECT 668.870 1577.130 671.770 1577.190 ;
        RECT 848.870 1577.130 851.770 1577.190 ;
        RECT 1028.870 1577.130 1031.770 1577.190 ;
        RECT 1208.870 1577.130 1211.770 1577.190 ;
        RECT 1388.870 1577.130 1391.770 1577.190 ;
        RECT 1568.870 1577.130 1571.770 1577.190 ;
        RECT 1748.870 1577.130 1751.770 1577.190 ;
        RECT 1928.870 1577.130 1931.770 1577.190 ;
        RECT 2108.870 1577.130 2111.770 1577.190 ;
        RECT 2288.870 1577.130 2291.770 1577.190 ;
        RECT 2468.870 1577.130 2471.770 1577.190 ;
        RECT 2648.870 1577.130 2651.770 1577.190 ;
        RECT 2828.870 1577.130 2831.770 1577.190 ;
        RECT 2949.650 1577.130 2952.550 1577.190 ;
        RECT -32.930 1574.230 2952.550 1577.130 ;
        RECT -32.930 1574.170 -30.030 1574.230 ;
        RECT 128.870 1574.170 131.770 1574.230 ;
        RECT 308.870 1574.170 311.770 1574.230 ;
        RECT 488.870 1574.170 491.770 1574.230 ;
        RECT 668.870 1574.170 671.770 1574.230 ;
        RECT 848.870 1574.170 851.770 1574.230 ;
        RECT 1028.870 1574.170 1031.770 1574.230 ;
        RECT 1208.870 1574.170 1211.770 1574.230 ;
        RECT 1388.870 1574.170 1391.770 1574.230 ;
        RECT 1568.870 1574.170 1571.770 1574.230 ;
        RECT 1748.870 1574.170 1751.770 1574.230 ;
        RECT 1928.870 1574.170 1931.770 1574.230 ;
        RECT 2108.870 1574.170 2111.770 1574.230 ;
        RECT 2288.870 1574.170 2291.770 1574.230 ;
        RECT 2468.870 1574.170 2471.770 1574.230 ;
        RECT 2648.870 1574.170 2651.770 1574.230 ;
        RECT 2828.870 1574.170 2831.770 1574.230 ;
        RECT 2949.650 1574.170 2952.550 1574.230 ;
        RECT -32.930 1397.130 -30.030 1397.190 ;
        RECT 128.870 1397.130 131.770 1397.190 ;
        RECT 308.870 1397.130 311.770 1397.190 ;
        RECT 488.870 1397.130 491.770 1397.190 ;
        RECT 668.870 1397.130 671.770 1397.190 ;
        RECT 848.870 1397.130 851.770 1397.190 ;
        RECT 1028.870 1397.130 1031.770 1397.190 ;
        RECT 1208.870 1397.130 1211.770 1397.190 ;
        RECT 1388.870 1397.130 1391.770 1397.190 ;
        RECT 1568.870 1397.130 1571.770 1397.190 ;
        RECT 1748.870 1397.130 1751.770 1397.190 ;
        RECT 1928.870 1397.130 1931.770 1397.190 ;
        RECT 2108.870 1397.130 2111.770 1397.190 ;
        RECT 2288.870 1397.130 2291.770 1397.190 ;
        RECT 2468.870 1397.130 2471.770 1397.190 ;
        RECT 2648.870 1397.130 2651.770 1397.190 ;
        RECT 2828.870 1397.130 2831.770 1397.190 ;
        RECT 2949.650 1397.130 2952.550 1397.190 ;
        RECT -32.930 1394.230 2952.550 1397.130 ;
        RECT -32.930 1394.170 -30.030 1394.230 ;
        RECT 128.870 1394.170 131.770 1394.230 ;
        RECT 308.870 1394.170 311.770 1394.230 ;
        RECT 488.870 1394.170 491.770 1394.230 ;
        RECT 668.870 1394.170 671.770 1394.230 ;
        RECT 848.870 1394.170 851.770 1394.230 ;
        RECT 1028.870 1394.170 1031.770 1394.230 ;
        RECT 1208.870 1394.170 1211.770 1394.230 ;
        RECT 1388.870 1394.170 1391.770 1394.230 ;
        RECT 1568.870 1394.170 1571.770 1394.230 ;
        RECT 1748.870 1394.170 1751.770 1394.230 ;
        RECT 1928.870 1394.170 1931.770 1394.230 ;
        RECT 2108.870 1394.170 2111.770 1394.230 ;
        RECT 2288.870 1394.170 2291.770 1394.230 ;
        RECT 2468.870 1394.170 2471.770 1394.230 ;
        RECT 2648.870 1394.170 2651.770 1394.230 ;
        RECT 2828.870 1394.170 2831.770 1394.230 ;
        RECT 2949.650 1394.170 2952.550 1394.230 ;
        RECT -32.930 1217.130 -30.030 1217.190 ;
        RECT 128.870 1217.130 131.770 1217.190 ;
        RECT 308.870 1217.130 311.770 1217.190 ;
        RECT 488.870 1217.130 491.770 1217.190 ;
        RECT 668.870 1217.130 671.770 1217.190 ;
        RECT 848.870 1217.130 851.770 1217.190 ;
        RECT 1028.870 1217.130 1031.770 1217.190 ;
        RECT 1208.870 1217.130 1211.770 1217.190 ;
        RECT 1388.870 1217.130 1391.770 1217.190 ;
        RECT 1568.870 1217.130 1571.770 1217.190 ;
        RECT 1748.870 1217.130 1751.770 1217.190 ;
        RECT 1928.870 1217.130 1931.770 1217.190 ;
        RECT 2108.870 1217.130 2111.770 1217.190 ;
        RECT 2288.870 1217.130 2291.770 1217.190 ;
        RECT 2468.870 1217.130 2471.770 1217.190 ;
        RECT 2648.870 1217.130 2651.770 1217.190 ;
        RECT 2828.870 1217.130 2831.770 1217.190 ;
        RECT 2949.650 1217.130 2952.550 1217.190 ;
        RECT -32.930 1214.230 2952.550 1217.130 ;
        RECT -32.930 1214.170 -30.030 1214.230 ;
        RECT 128.870 1214.170 131.770 1214.230 ;
        RECT 308.870 1214.170 311.770 1214.230 ;
        RECT 488.870 1214.170 491.770 1214.230 ;
        RECT 668.870 1214.170 671.770 1214.230 ;
        RECT 848.870 1214.170 851.770 1214.230 ;
        RECT 1028.870 1214.170 1031.770 1214.230 ;
        RECT 1208.870 1214.170 1211.770 1214.230 ;
        RECT 1388.870 1214.170 1391.770 1214.230 ;
        RECT 1568.870 1214.170 1571.770 1214.230 ;
        RECT 1748.870 1214.170 1751.770 1214.230 ;
        RECT 1928.870 1214.170 1931.770 1214.230 ;
        RECT 2108.870 1214.170 2111.770 1214.230 ;
        RECT 2288.870 1214.170 2291.770 1214.230 ;
        RECT 2468.870 1214.170 2471.770 1214.230 ;
        RECT 2648.870 1214.170 2651.770 1214.230 ;
        RECT 2828.870 1214.170 2831.770 1214.230 ;
        RECT 2949.650 1214.170 2952.550 1214.230 ;
        RECT -32.930 1037.130 -30.030 1037.190 ;
        RECT 128.870 1037.130 131.770 1037.190 ;
        RECT 308.870 1037.130 311.770 1037.190 ;
        RECT 488.870 1037.130 491.770 1037.190 ;
        RECT 668.870 1037.130 671.770 1037.190 ;
        RECT 848.870 1037.130 851.770 1037.190 ;
        RECT 1028.870 1037.130 1031.770 1037.190 ;
        RECT 1208.870 1037.130 1211.770 1037.190 ;
        RECT 1388.870 1037.130 1391.770 1037.190 ;
        RECT 1568.870 1037.130 1571.770 1037.190 ;
        RECT 1748.870 1037.130 1751.770 1037.190 ;
        RECT 1928.870 1037.130 1931.770 1037.190 ;
        RECT 2108.870 1037.130 2111.770 1037.190 ;
        RECT 2288.870 1037.130 2291.770 1037.190 ;
        RECT 2468.870 1037.130 2471.770 1037.190 ;
        RECT 2648.870 1037.130 2651.770 1037.190 ;
        RECT 2828.870 1037.130 2831.770 1037.190 ;
        RECT 2949.650 1037.130 2952.550 1037.190 ;
        RECT -32.930 1034.230 2952.550 1037.130 ;
        RECT -32.930 1034.170 -30.030 1034.230 ;
        RECT 128.870 1034.170 131.770 1034.230 ;
        RECT 308.870 1034.170 311.770 1034.230 ;
        RECT 488.870 1034.170 491.770 1034.230 ;
        RECT 668.870 1034.170 671.770 1034.230 ;
        RECT 848.870 1034.170 851.770 1034.230 ;
        RECT 1028.870 1034.170 1031.770 1034.230 ;
        RECT 1208.870 1034.170 1211.770 1034.230 ;
        RECT 1388.870 1034.170 1391.770 1034.230 ;
        RECT 1568.870 1034.170 1571.770 1034.230 ;
        RECT 1748.870 1034.170 1751.770 1034.230 ;
        RECT 1928.870 1034.170 1931.770 1034.230 ;
        RECT 2108.870 1034.170 2111.770 1034.230 ;
        RECT 2288.870 1034.170 2291.770 1034.230 ;
        RECT 2468.870 1034.170 2471.770 1034.230 ;
        RECT 2648.870 1034.170 2651.770 1034.230 ;
        RECT 2828.870 1034.170 2831.770 1034.230 ;
        RECT 2949.650 1034.170 2952.550 1034.230 ;
        RECT -32.930 857.130 -30.030 857.190 ;
        RECT 128.870 857.130 131.770 857.190 ;
        RECT 308.870 857.130 311.770 857.190 ;
        RECT 488.870 857.130 491.770 857.190 ;
        RECT 668.870 857.130 671.770 857.190 ;
        RECT 848.870 857.130 851.770 857.190 ;
        RECT 1028.870 857.130 1031.770 857.190 ;
        RECT 1208.870 857.130 1211.770 857.190 ;
        RECT 1388.870 857.130 1391.770 857.190 ;
        RECT 1568.870 857.130 1571.770 857.190 ;
        RECT 1748.870 857.130 1751.770 857.190 ;
        RECT 1928.870 857.130 1931.770 857.190 ;
        RECT 2108.870 857.130 2111.770 857.190 ;
        RECT 2288.870 857.130 2291.770 857.190 ;
        RECT 2468.870 857.130 2471.770 857.190 ;
        RECT 2648.870 857.130 2651.770 857.190 ;
        RECT 2828.870 857.130 2831.770 857.190 ;
        RECT 2949.650 857.130 2952.550 857.190 ;
        RECT -32.930 854.230 2952.550 857.130 ;
        RECT -32.930 854.170 -30.030 854.230 ;
        RECT 128.870 854.170 131.770 854.230 ;
        RECT 308.870 854.170 311.770 854.230 ;
        RECT 488.870 854.170 491.770 854.230 ;
        RECT 668.870 854.170 671.770 854.230 ;
        RECT 848.870 854.170 851.770 854.230 ;
        RECT 1028.870 854.170 1031.770 854.230 ;
        RECT 1208.870 854.170 1211.770 854.230 ;
        RECT 1388.870 854.170 1391.770 854.230 ;
        RECT 1568.870 854.170 1571.770 854.230 ;
        RECT 1748.870 854.170 1751.770 854.230 ;
        RECT 1928.870 854.170 1931.770 854.230 ;
        RECT 2108.870 854.170 2111.770 854.230 ;
        RECT 2288.870 854.170 2291.770 854.230 ;
        RECT 2468.870 854.170 2471.770 854.230 ;
        RECT 2648.870 854.170 2651.770 854.230 ;
        RECT 2828.870 854.170 2831.770 854.230 ;
        RECT 2949.650 854.170 2952.550 854.230 ;
        RECT -32.930 677.130 -30.030 677.190 ;
        RECT 128.870 677.130 131.770 677.190 ;
        RECT 308.870 677.130 311.770 677.190 ;
        RECT 488.870 677.130 491.770 677.190 ;
        RECT 668.870 677.130 671.770 677.190 ;
        RECT 848.870 677.130 851.770 677.190 ;
        RECT 1028.870 677.130 1031.770 677.190 ;
        RECT 1208.870 677.130 1211.770 677.190 ;
        RECT 1388.870 677.130 1391.770 677.190 ;
        RECT 1568.870 677.130 1571.770 677.190 ;
        RECT 1748.870 677.130 1751.770 677.190 ;
        RECT 1928.870 677.130 1931.770 677.190 ;
        RECT 2108.870 677.130 2111.770 677.190 ;
        RECT 2288.870 677.130 2291.770 677.190 ;
        RECT 2468.870 677.130 2471.770 677.190 ;
        RECT 2648.870 677.130 2651.770 677.190 ;
        RECT 2828.870 677.130 2831.770 677.190 ;
        RECT 2949.650 677.130 2952.550 677.190 ;
        RECT -32.930 674.230 2952.550 677.130 ;
        RECT -32.930 674.170 -30.030 674.230 ;
        RECT 128.870 674.170 131.770 674.230 ;
        RECT 308.870 674.170 311.770 674.230 ;
        RECT 488.870 674.170 491.770 674.230 ;
        RECT 668.870 674.170 671.770 674.230 ;
        RECT 848.870 674.170 851.770 674.230 ;
        RECT 1028.870 674.170 1031.770 674.230 ;
        RECT 1208.870 674.170 1211.770 674.230 ;
        RECT 1388.870 674.170 1391.770 674.230 ;
        RECT 1568.870 674.170 1571.770 674.230 ;
        RECT 1748.870 674.170 1751.770 674.230 ;
        RECT 1928.870 674.170 1931.770 674.230 ;
        RECT 2108.870 674.170 2111.770 674.230 ;
        RECT 2288.870 674.170 2291.770 674.230 ;
        RECT 2468.870 674.170 2471.770 674.230 ;
        RECT 2648.870 674.170 2651.770 674.230 ;
        RECT 2828.870 674.170 2831.770 674.230 ;
        RECT 2949.650 674.170 2952.550 674.230 ;
        RECT -32.930 497.130 -30.030 497.190 ;
        RECT 128.870 497.130 131.770 497.190 ;
        RECT 308.870 497.130 311.770 497.190 ;
        RECT 488.870 497.130 491.770 497.190 ;
        RECT 668.870 497.130 671.770 497.190 ;
        RECT 848.870 497.130 851.770 497.190 ;
        RECT 1028.870 497.130 1031.770 497.190 ;
        RECT 1208.870 497.130 1211.770 497.190 ;
        RECT 1388.870 497.130 1391.770 497.190 ;
        RECT 1568.870 497.130 1571.770 497.190 ;
        RECT 1748.870 497.130 1751.770 497.190 ;
        RECT 1928.870 497.130 1931.770 497.190 ;
        RECT 2108.870 497.130 2111.770 497.190 ;
        RECT 2288.870 497.130 2291.770 497.190 ;
        RECT 2468.870 497.130 2471.770 497.190 ;
        RECT 2648.870 497.130 2651.770 497.190 ;
        RECT 2828.870 497.130 2831.770 497.190 ;
        RECT 2949.650 497.130 2952.550 497.190 ;
        RECT -32.930 494.230 2952.550 497.130 ;
        RECT -32.930 494.170 -30.030 494.230 ;
        RECT 128.870 494.170 131.770 494.230 ;
        RECT 308.870 494.170 311.770 494.230 ;
        RECT 488.870 494.170 491.770 494.230 ;
        RECT 668.870 494.170 671.770 494.230 ;
        RECT 848.870 494.170 851.770 494.230 ;
        RECT 1028.870 494.170 1031.770 494.230 ;
        RECT 1208.870 494.170 1211.770 494.230 ;
        RECT 1388.870 494.170 1391.770 494.230 ;
        RECT 1568.870 494.170 1571.770 494.230 ;
        RECT 1748.870 494.170 1751.770 494.230 ;
        RECT 1928.870 494.170 1931.770 494.230 ;
        RECT 2108.870 494.170 2111.770 494.230 ;
        RECT 2288.870 494.170 2291.770 494.230 ;
        RECT 2468.870 494.170 2471.770 494.230 ;
        RECT 2648.870 494.170 2651.770 494.230 ;
        RECT 2828.870 494.170 2831.770 494.230 ;
        RECT 2949.650 494.170 2952.550 494.230 ;
        RECT -32.930 317.130 -30.030 317.190 ;
        RECT 128.870 317.130 131.770 317.190 ;
        RECT 308.870 317.130 311.770 317.190 ;
        RECT 488.870 317.130 491.770 317.190 ;
        RECT 668.870 317.130 671.770 317.190 ;
        RECT 848.870 317.130 851.770 317.190 ;
        RECT 1028.870 317.130 1031.770 317.190 ;
        RECT 1208.870 317.130 1211.770 317.190 ;
        RECT 1388.870 317.130 1391.770 317.190 ;
        RECT 1568.870 317.130 1571.770 317.190 ;
        RECT 1748.870 317.130 1751.770 317.190 ;
        RECT 1928.870 317.130 1931.770 317.190 ;
        RECT 2108.870 317.130 2111.770 317.190 ;
        RECT 2288.870 317.130 2291.770 317.190 ;
        RECT 2468.870 317.130 2471.770 317.190 ;
        RECT 2648.870 317.130 2651.770 317.190 ;
        RECT 2828.870 317.130 2831.770 317.190 ;
        RECT 2949.650 317.130 2952.550 317.190 ;
        RECT -32.930 314.230 2952.550 317.130 ;
        RECT -32.930 314.170 -30.030 314.230 ;
        RECT 128.870 314.170 131.770 314.230 ;
        RECT 308.870 314.170 311.770 314.230 ;
        RECT 488.870 314.170 491.770 314.230 ;
        RECT 668.870 314.170 671.770 314.230 ;
        RECT 848.870 314.170 851.770 314.230 ;
        RECT 1028.870 314.170 1031.770 314.230 ;
        RECT 1208.870 314.170 1211.770 314.230 ;
        RECT 1388.870 314.170 1391.770 314.230 ;
        RECT 1568.870 314.170 1571.770 314.230 ;
        RECT 1748.870 314.170 1751.770 314.230 ;
        RECT 1928.870 314.170 1931.770 314.230 ;
        RECT 2108.870 314.170 2111.770 314.230 ;
        RECT 2288.870 314.170 2291.770 314.230 ;
        RECT 2468.870 314.170 2471.770 314.230 ;
        RECT 2648.870 314.170 2651.770 314.230 ;
        RECT 2828.870 314.170 2831.770 314.230 ;
        RECT 2949.650 314.170 2952.550 314.230 ;
        RECT -32.930 137.130 -30.030 137.190 ;
        RECT 128.870 137.130 131.770 137.190 ;
        RECT 308.870 137.130 311.770 137.190 ;
        RECT 488.870 137.130 491.770 137.190 ;
        RECT 668.870 137.130 671.770 137.190 ;
        RECT 848.870 137.130 851.770 137.190 ;
        RECT 1028.870 137.130 1031.770 137.190 ;
        RECT 1208.870 137.130 1211.770 137.190 ;
        RECT 1388.870 137.130 1391.770 137.190 ;
        RECT 1568.870 137.130 1571.770 137.190 ;
        RECT 1748.870 137.130 1751.770 137.190 ;
        RECT 1928.870 137.130 1931.770 137.190 ;
        RECT 2108.870 137.130 2111.770 137.190 ;
        RECT 2288.870 137.130 2291.770 137.190 ;
        RECT 2468.870 137.130 2471.770 137.190 ;
        RECT 2648.870 137.130 2651.770 137.190 ;
        RECT 2828.870 137.130 2831.770 137.190 ;
        RECT 2949.650 137.130 2952.550 137.190 ;
        RECT -32.930 134.230 2952.550 137.130 ;
        RECT -32.930 134.170 -30.030 134.230 ;
        RECT 128.870 134.170 131.770 134.230 ;
        RECT 308.870 134.170 311.770 134.230 ;
        RECT 488.870 134.170 491.770 134.230 ;
        RECT 668.870 134.170 671.770 134.230 ;
        RECT 848.870 134.170 851.770 134.230 ;
        RECT 1028.870 134.170 1031.770 134.230 ;
        RECT 1208.870 134.170 1211.770 134.230 ;
        RECT 1388.870 134.170 1391.770 134.230 ;
        RECT 1568.870 134.170 1571.770 134.230 ;
        RECT 1748.870 134.170 1751.770 134.230 ;
        RECT 1928.870 134.170 1931.770 134.230 ;
        RECT 2108.870 134.170 2111.770 134.230 ;
        RECT 2288.870 134.170 2291.770 134.230 ;
        RECT 2468.870 134.170 2471.770 134.230 ;
        RECT 2648.870 134.170 2651.770 134.230 ;
        RECT 2828.870 134.170 2831.770 134.230 ;
        RECT 2949.650 134.170 2952.550 134.230 ;
        RECT -32.930 -24.670 -30.030 -24.610 ;
        RECT 128.870 -24.670 131.770 -24.610 ;
        RECT 308.870 -24.670 311.770 -24.610 ;
        RECT 488.870 -24.670 491.770 -24.610 ;
        RECT 668.870 -24.670 671.770 -24.610 ;
        RECT 848.870 -24.670 851.770 -24.610 ;
        RECT 1028.870 -24.670 1031.770 -24.610 ;
        RECT 1208.870 -24.670 1211.770 -24.610 ;
        RECT 1388.870 -24.670 1391.770 -24.610 ;
        RECT 1568.870 -24.670 1571.770 -24.610 ;
        RECT 1748.870 -24.670 1751.770 -24.610 ;
        RECT 1928.870 -24.670 1931.770 -24.610 ;
        RECT 2108.870 -24.670 2111.770 -24.610 ;
        RECT 2288.870 -24.670 2291.770 -24.610 ;
        RECT 2468.870 -24.670 2471.770 -24.610 ;
        RECT 2648.870 -24.670 2651.770 -24.610 ;
        RECT 2828.870 -24.670 2831.770 -24.610 ;
        RECT 2949.650 -24.670 2952.550 -24.610 ;
        RECT -32.930 -27.570 2952.550 -24.670 ;
        RECT -32.930 -27.630 -30.030 -27.570 ;
        RECT 128.870 -27.630 131.770 -27.570 ;
        RECT 308.870 -27.630 311.770 -27.570 ;
        RECT 488.870 -27.630 491.770 -27.570 ;
        RECT 668.870 -27.630 671.770 -27.570 ;
        RECT 848.870 -27.630 851.770 -27.570 ;
        RECT 1028.870 -27.630 1031.770 -27.570 ;
        RECT 1208.870 -27.630 1211.770 -27.570 ;
        RECT 1388.870 -27.630 1391.770 -27.570 ;
        RECT 1568.870 -27.630 1571.770 -27.570 ;
        RECT 1748.870 -27.630 1751.770 -27.570 ;
        RECT 1928.870 -27.630 1931.770 -27.570 ;
        RECT 2108.870 -27.630 2111.770 -27.570 ;
        RECT 2288.870 -27.630 2291.770 -27.570 ;
        RECT 2468.870 -27.630 2471.770 -27.570 ;
        RECT 2648.870 -27.630 2651.770 -27.570 ;
        RECT 2828.870 -27.630 2831.770 -27.570 ;
        RECT 2949.650 -27.630 2952.550 -27.570 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.530 -32.170 -34.630 3551.850 ;
        RECT 56.270 -36.770 59.170 3556.450 ;
        RECT 236.270 -36.770 239.170 3556.450 ;
        RECT 416.270 -36.770 419.170 3556.450 ;
        RECT 596.270 -36.770 599.170 3556.450 ;
        RECT 776.270 -36.770 779.170 3556.450 ;
        RECT 956.270 -36.770 959.170 3556.450 ;
        RECT 1136.270 -36.770 1139.170 3556.450 ;
        RECT 1316.270 -36.770 1319.170 3556.450 ;
        RECT 1496.270 -36.770 1499.170 3556.450 ;
        RECT 1676.270 -36.770 1679.170 3556.450 ;
        RECT 1856.270 -36.770 1859.170 3556.450 ;
        RECT 2036.270 -36.770 2039.170 3556.450 ;
        RECT 2216.270 -36.770 2219.170 3556.450 ;
        RECT 2396.270 -36.770 2399.170 3556.450 ;
        RECT 2576.270 -36.770 2579.170 3556.450 ;
        RECT 2756.270 -36.770 2759.170 3556.450 ;
        RECT 2954.250 -32.170 2957.150 3551.850 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3483.290 -35.490 3484.470 ;
        RECT -36.670 3481.690 -35.490 3482.870 ;
        RECT -36.670 3303.290 -35.490 3304.470 ;
        RECT -36.670 3301.690 -35.490 3302.870 ;
        RECT -36.670 3123.290 -35.490 3124.470 ;
        RECT -36.670 3121.690 -35.490 3122.870 ;
        RECT -36.670 2943.290 -35.490 2944.470 ;
        RECT -36.670 2941.690 -35.490 2942.870 ;
        RECT -36.670 2763.290 -35.490 2764.470 ;
        RECT -36.670 2761.690 -35.490 2762.870 ;
        RECT -36.670 2583.290 -35.490 2584.470 ;
        RECT -36.670 2581.690 -35.490 2582.870 ;
        RECT -36.670 2403.290 -35.490 2404.470 ;
        RECT -36.670 2401.690 -35.490 2402.870 ;
        RECT -36.670 2223.290 -35.490 2224.470 ;
        RECT -36.670 2221.690 -35.490 2222.870 ;
        RECT -36.670 2043.290 -35.490 2044.470 ;
        RECT -36.670 2041.690 -35.490 2042.870 ;
        RECT -36.670 1863.290 -35.490 1864.470 ;
        RECT -36.670 1861.690 -35.490 1862.870 ;
        RECT -36.670 1683.290 -35.490 1684.470 ;
        RECT -36.670 1681.690 -35.490 1682.870 ;
        RECT -36.670 1503.290 -35.490 1504.470 ;
        RECT -36.670 1501.690 -35.490 1502.870 ;
        RECT -36.670 1323.290 -35.490 1324.470 ;
        RECT -36.670 1321.690 -35.490 1322.870 ;
        RECT -36.670 1143.290 -35.490 1144.470 ;
        RECT -36.670 1141.690 -35.490 1142.870 ;
        RECT -36.670 963.290 -35.490 964.470 ;
        RECT -36.670 961.690 -35.490 962.870 ;
        RECT -36.670 783.290 -35.490 784.470 ;
        RECT -36.670 781.690 -35.490 782.870 ;
        RECT -36.670 603.290 -35.490 604.470 ;
        RECT -36.670 601.690 -35.490 602.870 ;
        RECT -36.670 423.290 -35.490 424.470 ;
        RECT -36.670 421.690 -35.490 422.870 ;
        RECT -36.670 243.290 -35.490 244.470 ;
        RECT -36.670 241.690 -35.490 242.870 ;
        RECT -36.670 63.290 -35.490 64.470 ;
        RECT -36.670 61.690 -35.490 62.870 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 57.130 3550.610 58.310 3551.790 ;
        RECT 57.130 3549.010 58.310 3550.190 ;
        RECT 57.130 3483.290 58.310 3484.470 ;
        RECT 57.130 3481.690 58.310 3482.870 ;
        RECT 57.130 3303.290 58.310 3304.470 ;
        RECT 57.130 3301.690 58.310 3302.870 ;
        RECT 57.130 3123.290 58.310 3124.470 ;
        RECT 57.130 3121.690 58.310 3122.870 ;
        RECT 57.130 2943.290 58.310 2944.470 ;
        RECT 57.130 2941.690 58.310 2942.870 ;
        RECT 57.130 2763.290 58.310 2764.470 ;
        RECT 57.130 2761.690 58.310 2762.870 ;
        RECT 57.130 2583.290 58.310 2584.470 ;
        RECT 57.130 2581.690 58.310 2582.870 ;
        RECT 57.130 2403.290 58.310 2404.470 ;
        RECT 57.130 2401.690 58.310 2402.870 ;
        RECT 57.130 2223.290 58.310 2224.470 ;
        RECT 57.130 2221.690 58.310 2222.870 ;
        RECT 57.130 2043.290 58.310 2044.470 ;
        RECT 57.130 2041.690 58.310 2042.870 ;
        RECT 57.130 1863.290 58.310 1864.470 ;
        RECT 57.130 1861.690 58.310 1862.870 ;
        RECT 57.130 1683.290 58.310 1684.470 ;
        RECT 57.130 1681.690 58.310 1682.870 ;
        RECT 57.130 1503.290 58.310 1504.470 ;
        RECT 57.130 1501.690 58.310 1502.870 ;
        RECT 57.130 1323.290 58.310 1324.470 ;
        RECT 57.130 1321.690 58.310 1322.870 ;
        RECT 57.130 1143.290 58.310 1144.470 ;
        RECT 57.130 1141.690 58.310 1142.870 ;
        RECT 57.130 963.290 58.310 964.470 ;
        RECT 57.130 961.690 58.310 962.870 ;
        RECT 57.130 783.290 58.310 784.470 ;
        RECT 57.130 781.690 58.310 782.870 ;
        RECT 57.130 603.290 58.310 604.470 ;
        RECT 57.130 601.690 58.310 602.870 ;
        RECT 57.130 423.290 58.310 424.470 ;
        RECT 57.130 421.690 58.310 422.870 ;
        RECT 57.130 243.290 58.310 244.470 ;
        RECT 57.130 241.690 58.310 242.870 ;
        RECT 57.130 63.290 58.310 64.470 ;
        RECT 57.130 61.690 58.310 62.870 ;
        RECT 57.130 -30.510 58.310 -29.330 ;
        RECT 57.130 -32.110 58.310 -30.930 ;
        RECT 237.130 3550.610 238.310 3551.790 ;
        RECT 237.130 3549.010 238.310 3550.190 ;
        RECT 237.130 3483.290 238.310 3484.470 ;
        RECT 237.130 3481.690 238.310 3482.870 ;
        RECT 237.130 3303.290 238.310 3304.470 ;
        RECT 237.130 3301.690 238.310 3302.870 ;
        RECT 237.130 3123.290 238.310 3124.470 ;
        RECT 237.130 3121.690 238.310 3122.870 ;
        RECT 237.130 2943.290 238.310 2944.470 ;
        RECT 237.130 2941.690 238.310 2942.870 ;
        RECT 237.130 2763.290 238.310 2764.470 ;
        RECT 237.130 2761.690 238.310 2762.870 ;
        RECT 237.130 2583.290 238.310 2584.470 ;
        RECT 237.130 2581.690 238.310 2582.870 ;
        RECT 237.130 2403.290 238.310 2404.470 ;
        RECT 237.130 2401.690 238.310 2402.870 ;
        RECT 237.130 2223.290 238.310 2224.470 ;
        RECT 237.130 2221.690 238.310 2222.870 ;
        RECT 237.130 2043.290 238.310 2044.470 ;
        RECT 237.130 2041.690 238.310 2042.870 ;
        RECT 237.130 1863.290 238.310 1864.470 ;
        RECT 237.130 1861.690 238.310 1862.870 ;
        RECT 237.130 1683.290 238.310 1684.470 ;
        RECT 237.130 1681.690 238.310 1682.870 ;
        RECT 237.130 1503.290 238.310 1504.470 ;
        RECT 237.130 1501.690 238.310 1502.870 ;
        RECT 237.130 1323.290 238.310 1324.470 ;
        RECT 237.130 1321.690 238.310 1322.870 ;
        RECT 237.130 1143.290 238.310 1144.470 ;
        RECT 237.130 1141.690 238.310 1142.870 ;
        RECT 237.130 963.290 238.310 964.470 ;
        RECT 237.130 961.690 238.310 962.870 ;
        RECT 237.130 783.290 238.310 784.470 ;
        RECT 237.130 781.690 238.310 782.870 ;
        RECT 237.130 603.290 238.310 604.470 ;
        RECT 237.130 601.690 238.310 602.870 ;
        RECT 237.130 423.290 238.310 424.470 ;
        RECT 237.130 421.690 238.310 422.870 ;
        RECT 237.130 243.290 238.310 244.470 ;
        RECT 237.130 241.690 238.310 242.870 ;
        RECT 237.130 63.290 238.310 64.470 ;
        RECT 237.130 61.690 238.310 62.870 ;
        RECT 237.130 -30.510 238.310 -29.330 ;
        RECT 237.130 -32.110 238.310 -30.930 ;
        RECT 417.130 3550.610 418.310 3551.790 ;
        RECT 417.130 3549.010 418.310 3550.190 ;
        RECT 417.130 3483.290 418.310 3484.470 ;
        RECT 417.130 3481.690 418.310 3482.870 ;
        RECT 417.130 3303.290 418.310 3304.470 ;
        RECT 417.130 3301.690 418.310 3302.870 ;
        RECT 417.130 3123.290 418.310 3124.470 ;
        RECT 417.130 3121.690 418.310 3122.870 ;
        RECT 417.130 2943.290 418.310 2944.470 ;
        RECT 417.130 2941.690 418.310 2942.870 ;
        RECT 417.130 2763.290 418.310 2764.470 ;
        RECT 417.130 2761.690 418.310 2762.870 ;
        RECT 417.130 2583.290 418.310 2584.470 ;
        RECT 417.130 2581.690 418.310 2582.870 ;
        RECT 417.130 2403.290 418.310 2404.470 ;
        RECT 417.130 2401.690 418.310 2402.870 ;
        RECT 417.130 2223.290 418.310 2224.470 ;
        RECT 417.130 2221.690 418.310 2222.870 ;
        RECT 417.130 2043.290 418.310 2044.470 ;
        RECT 417.130 2041.690 418.310 2042.870 ;
        RECT 417.130 1863.290 418.310 1864.470 ;
        RECT 417.130 1861.690 418.310 1862.870 ;
        RECT 417.130 1683.290 418.310 1684.470 ;
        RECT 417.130 1681.690 418.310 1682.870 ;
        RECT 417.130 1503.290 418.310 1504.470 ;
        RECT 417.130 1501.690 418.310 1502.870 ;
        RECT 417.130 1323.290 418.310 1324.470 ;
        RECT 417.130 1321.690 418.310 1322.870 ;
        RECT 417.130 1143.290 418.310 1144.470 ;
        RECT 417.130 1141.690 418.310 1142.870 ;
        RECT 417.130 963.290 418.310 964.470 ;
        RECT 417.130 961.690 418.310 962.870 ;
        RECT 417.130 783.290 418.310 784.470 ;
        RECT 417.130 781.690 418.310 782.870 ;
        RECT 417.130 603.290 418.310 604.470 ;
        RECT 417.130 601.690 418.310 602.870 ;
        RECT 417.130 423.290 418.310 424.470 ;
        RECT 417.130 421.690 418.310 422.870 ;
        RECT 417.130 243.290 418.310 244.470 ;
        RECT 417.130 241.690 418.310 242.870 ;
        RECT 417.130 63.290 418.310 64.470 ;
        RECT 417.130 61.690 418.310 62.870 ;
        RECT 417.130 -30.510 418.310 -29.330 ;
        RECT 417.130 -32.110 418.310 -30.930 ;
        RECT 597.130 3550.610 598.310 3551.790 ;
        RECT 597.130 3549.010 598.310 3550.190 ;
        RECT 597.130 3483.290 598.310 3484.470 ;
        RECT 597.130 3481.690 598.310 3482.870 ;
        RECT 597.130 3303.290 598.310 3304.470 ;
        RECT 597.130 3301.690 598.310 3302.870 ;
        RECT 597.130 3123.290 598.310 3124.470 ;
        RECT 597.130 3121.690 598.310 3122.870 ;
        RECT 597.130 2943.290 598.310 2944.470 ;
        RECT 597.130 2941.690 598.310 2942.870 ;
        RECT 597.130 2763.290 598.310 2764.470 ;
        RECT 597.130 2761.690 598.310 2762.870 ;
        RECT 597.130 2583.290 598.310 2584.470 ;
        RECT 597.130 2581.690 598.310 2582.870 ;
        RECT 597.130 2403.290 598.310 2404.470 ;
        RECT 597.130 2401.690 598.310 2402.870 ;
        RECT 597.130 2223.290 598.310 2224.470 ;
        RECT 597.130 2221.690 598.310 2222.870 ;
        RECT 597.130 2043.290 598.310 2044.470 ;
        RECT 597.130 2041.690 598.310 2042.870 ;
        RECT 597.130 1863.290 598.310 1864.470 ;
        RECT 597.130 1861.690 598.310 1862.870 ;
        RECT 597.130 1683.290 598.310 1684.470 ;
        RECT 597.130 1681.690 598.310 1682.870 ;
        RECT 597.130 1503.290 598.310 1504.470 ;
        RECT 597.130 1501.690 598.310 1502.870 ;
        RECT 597.130 1323.290 598.310 1324.470 ;
        RECT 597.130 1321.690 598.310 1322.870 ;
        RECT 597.130 1143.290 598.310 1144.470 ;
        RECT 597.130 1141.690 598.310 1142.870 ;
        RECT 597.130 963.290 598.310 964.470 ;
        RECT 597.130 961.690 598.310 962.870 ;
        RECT 597.130 783.290 598.310 784.470 ;
        RECT 597.130 781.690 598.310 782.870 ;
        RECT 597.130 603.290 598.310 604.470 ;
        RECT 597.130 601.690 598.310 602.870 ;
        RECT 597.130 423.290 598.310 424.470 ;
        RECT 597.130 421.690 598.310 422.870 ;
        RECT 597.130 243.290 598.310 244.470 ;
        RECT 597.130 241.690 598.310 242.870 ;
        RECT 597.130 63.290 598.310 64.470 ;
        RECT 597.130 61.690 598.310 62.870 ;
        RECT 597.130 -30.510 598.310 -29.330 ;
        RECT 597.130 -32.110 598.310 -30.930 ;
        RECT 777.130 3550.610 778.310 3551.790 ;
        RECT 777.130 3549.010 778.310 3550.190 ;
        RECT 777.130 3483.290 778.310 3484.470 ;
        RECT 777.130 3481.690 778.310 3482.870 ;
        RECT 777.130 3303.290 778.310 3304.470 ;
        RECT 777.130 3301.690 778.310 3302.870 ;
        RECT 777.130 3123.290 778.310 3124.470 ;
        RECT 777.130 3121.690 778.310 3122.870 ;
        RECT 777.130 2943.290 778.310 2944.470 ;
        RECT 777.130 2941.690 778.310 2942.870 ;
        RECT 777.130 2763.290 778.310 2764.470 ;
        RECT 777.130 2761.690 778.310 2762.870 ;
        RECT 777.130 2583.290 778.310 2584.470 ;
        RECT 777.130 2581.690 778.310 2582.870 ;
        RECT 777.130 2403.290 778.310 2404.470 ;
        RECT 777.130 2401.690 778.310 2402.870 ;
        RECT 777.130 2223.290 778.310 2224.470 ;
        RECT 777.130 2221.690 778.310 2222.870 ;
        RECT 777.130 2043.290 778.310 2044.470 ;
        RECT 777.130 2041.690 778.310 2042.870 ;
        RECT 777.130 1863.290 778.310 1864.470 ;
        RECT 777.130 1861.690 778.310 1862.870 ;
        RECT 777.130 1683.290 778.310 1684.470 ;
        RECT 777.130 1681.690 778.310 1682.870 ;
        RECT 777.130 1503.290 778.310 1504.470 ;
        RECT 777.130 1501.690 778.310 1502.870 ;
        RECT 777.130 1323.290 778.310 1324.470 ;
        RECT 777.130 1321.690 778.310 1322.870 ;
        RECT 777.130 1143.290 778.310 1144.470 ;
        RECT 777.130 1141.690 778.310 1142.870 ;
        RECT 777.130 963.290 778.310 964.470 ;
        RECT 777.130 961.690 778.310 962.870 ;
        RECT 777.130 783.290 778.310 784.470 ;
        RECT 777.130 781.690 778.310 782.870 ;
        RECT 777.130 603.290 778.310 604.470 ;
        RECT 777.130 601.690 778.310 602.870 ;
        RECT 777.130 423.290 778.310 424.470 ;
        RECT 777.130 421.690 778.310 422.870 ;
        RECT 777.130 243.290 778.310 244.470 ;
        RECT 777.130 241.690 778.310 242.870 ;
        RECT 777.130 63.290 778.310 64.470 ;
        RECT 777.130 61.690 778.310 62.870 ;
        RECT 777.130 -30.510 778.310 -29.330 ;
        RECT 777.130 -32.110 778.310 -30.930 ;
        RECT 957.130 3550.610 958.310 3551.790 ;
        RECT 957.130 3549.010 958.310 3550.190 ;
        RECT 957.130 3483.290 958.310 3484.470 ;
        RECT 957.130 3481.690 958.310 3482.870 ;
        RECT 957.130 3303.290 958.310 3304.470 ;
        RECT 957.130 3301.690 958.310 3302.870 ;
        RECT 957.130 3123.290 958.310 3124.470 ;
        RECT 957.130 3121.690 958.310 3122.870 ;
        RECT 957.130 2943.290 958.310 2944.470 ;
        RECT 957.130 2941.690 958.310 2942.870 ;
        RECT 957.130 2763.290 958.310 2764.470 ;
        RECT 957.130 2761.690 958.310 2762.870 ;
        RECT 957.130 2583.290 958.310 2584.470 ;
        RECT 957.130 2581.690 958.310 2582.870 ;
        RECT 957.130 2403.290 958.310 2404.470 ;
        RECT 957.130 2401.690 958.310 2402.870 ;
        RECT 957.130 2223.290 958.310 2224.470 ;
        RECT 957.130 2221.690 958.310 2222.870 ;
        RECT 957.130 2043.290 958.310 2044.470 ;
        RECT 957.130 2041.690 958.310 2042.870 ;
        RECT 957.130 1863.290 958.310 1864.470 ;
        RECT 957.130 1861.690 958.310 1862.870 ;
        RECT 957.130 1683.290 958.310 1684.470 ;
        RECT 957.130 1681.690 958.310 1682.870 ;
        RECT 957.130 1503.290 958.310 1504.470 ;
        RECT 957.130 1501.690 958.310 1502.870 ;
        RECT 957.130 1323.290 958.310 1324.470 ;
        RECT 957.130 1321.690 958.310 1322.870 ;
        RECT 957.130 1143.290 958.310 1144.470 ;
        RECT 957.130 1141.690 958.310 1142.870 ;
        RECT 957.130 963.290 958.310 964.470 ;
        RECT 957.130 961.690 958.310 962.870 ;
        RECT 957.130 783.290 958.310 784.470 ;
        RECT 957.130 781.690 958.310 782.870 ;
        RECT 957.130 603.290 958.310 604.470 ;
        RECT 957.130 601.690 958.310 602.870 ;
        RECT 957.130 423.290 958.310 424.470 ;
        RECT 957.130 421.690 958.310 422.870 ;
        RECT 957.130 243.290 958.310 244.470 ;
        RECT 957.130 241.690 958.310 242.870 ;
        RECT 957.130 63.290 958.310 64.470 ;
        RECT 957.130 61.690 958.310 62.870 ;
        RECT 957.130 -30.510 958.310 -29.330 ;
        RECT 957.130 -32.110 958.310 -30.930 ;
        RECT 1137.130 3550.610 1138.310 3551.790 ;
        RECT 1137.130 3549.010 1138.310 3550.190 ;
        RECT 1137.130 3483.290 1138.310 3484.470 ;
        RECT 1137.130 3481.690 1138.310 3482.870 ;
        RECT 1137.130 3303.290 1138.310 3304.470 ;
        RECT 1137.130 3301.690 1138.310 3302.870 ;
        RECT 1137.130 3123.290 1138.310 3124.470 ;
        RECT 1137.130 3121.690 1138.310 3122.870 ;
        RECT 1137.130 2943.290 1138.310 2944.470 ;
        RECT 1137.130 2941.690 1138.310 2942.870 ;
        RECT 1137.130 2763.290 1138.310 2764.470 ;
        RECT 1137.130 2761.690 1138.310 2762.870 ;
        RECT 1137.130 2583.290 1138.310 2584.470 ;
        RECT 1137.130 2581.690 1138.310 2582.870 ;
        RECT 1137.130 2403.290 1138.310 2404.470 ;
        RECT 1137.130 2401.690 1138.310 2402.870 ;
        RECT 1137.130 2223.290 1138.310 2224.470 ;
        RECT 1137.130 2221.690 1138.310 2222.870 ;
        RECT 1137.130 2043.290 1138.310 2044.470 ;
        RECT 1137.130 2041.690 1138.310 2042.870 ;
        RECT 1137.130 1863.290 1138.310 1864.470 ;
        RECT 1137.130 1861.690 1138.310 1862.870 ;
        RECT 1137.130 1683.290 1138.310 1684.470 ;
        RECT 1137.130 1681.690 1138.310 1682.870 ;
        RECT 1137.130 1503.290 1138.310 1504.470 ;
        RECT 1137.130 1501.690 1138.310 1502.870 ;
        RECT 1137.130 1323.290 1138.310 1324.470 ;
        RECT 1137.130 1321.690 1138.310 1322.870 ;
        RECT 1137.130 1143.290 1138.310 1144.470 ;
        RECT 1137.130 1141.690 1138.310 1142.870 ;
        RECT 1137.130 963.290 1138.310 964.470 ;
        RECT 1137.130 961.690 1138.310 962.870 ;
        RECT 1137.130 783.290 1138.310 784.470 ;
        RECT 1137.130 781.690 1138.310 782.870 ;
        RECT 1137.130 603.290 1138.310 604.470 ;
        RECT 1137.130 601.690 1138.310 602.870 ;
        RECT 1137.130 423.290 1138.310 424.470 ;
        RECT 1137.130 421.690 1138.310 422.870 ;
        RECT 1137.130 243.290 1138.310 244.470 ;
        RECT 1137.130 241.690 1138.310 242.870 ;
        RECT 1137.130 63.290 1138.310 64.470 ;
        RECT 1137.130 61.690 1138.310 62.870 ;
        RECT 1137.130 -30.510 1138.310 -29.330 ;
        RECT 1137.130 -32.110 1138.310 -30.930 ;
        RECT 1317.130 3550.610 1318.310 3551.790 ;
        RECT 1317.130 3549.010 1318.310 3550.190 ;
        RECT 1317.130 3483.290 1318.310 3484.470 ;
        RECT 1317.130 3481.690 1318.310 3482.870 ;
        RECT 1317.130 3303.290 1318.310 3304.470 ;
        RECT 1317.130 3301.690 1318.310 3302.870 ;
        RECT 1317.130 3123.290 1318.310 3124.470 ;
        RECT 1317.130 3121.690 1318.310 3122.870 ;
        RECT 1317.130 2943.290 1318.310 2944.470 ;
        RECT 1317.130 2941.690 1318.310 2942.870 ;
        RECT 1317.130 2763.290 1318.310 2764.470 ;
        RECT 1317.130 2761.690 1318.310 2762.870 ;
        RECT 1317.130 2583.290 1318.310 2584.470 ;
        RECT 1317.130 2581.690 1318.310 2582.870 ;
        RECT 1317.130 2403.290 1318.310 2404.470 ;
        RECT 1317.130 2401.690 1318.310 2402.870 ;
        RECT 1317.130 2223.290 1318.310 2224.470 ;
        RECT 1317.130 2221.690 1318.310 2222.870 ;
        RECT 1317.130 2043.290 1318.310 2044.470 ;
        RECT 1317.130 2041.690 1318.310 2042.870 ;
        RECT 1317.130 1863.290 1318.310 1864.470 ;
        RECT 1317.130 1861.690 1318.310 1862.870 ;
        RECT 1317.130 1683.290 1318.310 1684.470 ;
        RECT 1317.130 1681.690 1318.310 1682.870 ;
        RECT 1317.130 1503.290 1318.310 1504.470 ;
        RECT 1317.130 1501.690 1318.310 1502.870 ;
        RECT 1317.130 1323.290 1318.310 1324.470 ;
        RECT 1317.130 1321.690 1318.310 1322.870 ;
        RECT 1317.130 1143.290 1318.310 1144.470 ;
        RECT 1317.130 1141.690 1318.310 1142.870 ;
        RECT 1317.130 963.290 1318.310 964.470 ;
        RECT 1317.130 961.690 1318.310 962.870 ;
        RECT 1317.130 783.290 1318.310 784.470 ;
        RECT 1317.130 781.690 1318.310 782.870 ;
        RECT 1317.130 603.290 1318.310 604.470 ;
        RECT 1317.130 601.690 1318.310 602.870 ;
        RECT 1317.130 423.290 1318.310 424.470 ;
        RECT 1317.130 421.690 1318.310 422.870 ;
        RECT 1317.130 243.290 1318.310 244.470 ;
        RECT 1317.130 241.690 1318.310 242.870 ;
        RECT 1317.130 63.290 1318.310 64.470 ;
        RECT 1317.130 61.690 1318.310 62.870 ;
        RECT 1317.130 -30.510 1318.310 -29.330 ;
        RECT 1317.130 -32.110 1318.310 -30.930 ;
        RECT 1497.130 3550.610 1498.310 3551.790 ;
        RECT 1497.130 3549.010 1498.310 3550.190 ;
        RECT 1497.130 3483.290 1498.310 3484.470 ;
        RECT 1497.130 3481.690 1498.310 3482.870 ;
        RECT 1497.130 3303.290 1498.310 3304.470 ;
        RECT 1497.130 3301.690 1498.310 3302.870 ;
        RECT 1497.130 3123.290 1498.310 3124.470 ;
        RECT 1497.130 3121.690 1498.310 3122.870 ;
        RECT 1497.130 2943.290 1498.310 2944.470 ;
        RECT 1497.130 2941.690 1498.310 2942.870 ;
        RECT 1497.130 2763.290 1498.310 2764.470 ;
        RECT 1497.130 2761.690 1498.310 2762.870 ;
        RECT 1497.130 2583.290 1498.310 2584.470 ;
        RECT 1497.130 2581.690 1498.310 2582.870 ;
        RECT 1497.130 2403.290 1498.310 2404.470 ;
        RECT 1497.130 2401.690 1498.310 2402.870 ;
        RECT 1497.130 2223.290 1498.310 2224.470 ;
        RECT 1497.130 2221.690 1498.310 2222.870 ;
        RECT 1497.130 2043.290 1498.310 2044.470 ;
        RECT 1497.130 2041.690 1498.310 2042.870 ;
        RECT 1497.130 1863.290 1498.310 1864.470 ;
        RECT 1497.130 1861.690 1498.310 1862.870 ;
        RECT 1497.130 1683.290 1498.310 1684.470 ;
        RECT 1497.130 1681.690 1498.310 1682.870 ;
        RECT 1497.130 1503.290 1498.310 1504.470 ;
        RECT 1497.130 1501.690 1498.310 1502.870 ;
        RECT 1497.130 1323.290 1498.310 1324.470 ;
        RECT 1497.130 1321.690 1498.310 1322.870 ;
        RECT 1497.130 1143.290 1498.310 1144.470 ;
        RECT 1497.130 1141.690 1498.310 1142.870 ;
        RECT 1497.130 963.290 1498.310 964.470 ;
        RECT 1497.130 961.690 1498.310 962.870 ;
        RECT 1497.130 783.290 1498.310 784.470 ;
        RECT 1497.130 781.690 1498.310 782.870 ;
        RECT 1497.130 603.290 1498.310 604.470 ;
        RECT 1497.130 601.690 1498.310 602.870 ;
        RECT 1497.130 423.290 1498.310 424.470 ;
        RECT 1497.130 421.690 1498.310 422.870 ;
        RECT 1497.130 243.290 1498.310 244.470 ;
        RECT 1497.130 241.690 1498.310 242.870 ;
        RECT 1497.130 63.290 1498.310 64.470 ;
        RECT 1497.130 61.690 1498.310 62.870 ;
        RECT 1497.130 -30.510 1498.310 -29.330 ;
        RECT 1497.130 -32.110 1498.310 -30.930 ;
        RECT 1677.130 3550.610 1678.310 3551.790 ;
        RECT 1677.130 3549.010 1678.310 3550.190 ;
        RECT 1677.130 3483.290 1678.310 3484.470 ;
        RECT 1677.130 3481.690 1678.310 3482.870 ;
        RECT 1677.130 3303.290 1678.310 3304.470 ;
        RECT 1677.130 3301.690 1678.310 3302.870 ;
        RECT 1677.130 3123.290 1678.310 3124.470 ;
        RECT 1677.130 3121.690 1678.310 3122.870 ;
        RECT 1677.130 2943.290 1678.310 2944.470 ;
        RECT 1677.130 2941.690 1678.310 2942.870 ;
        RECT 1677.130 2763.290 1678.310 2764.470 ;
        RECT 1677.130 2761.690 1678.310 2762.870 ;
        RECT 1677.130 2583.290 1678.310 2584.470 ;
        RECT 1677.130 2581.690 1678.310 2582.870 ;
        RECT 1677.130 2403.290 1678.310 2404.470 ;
        RECT 1677.130 2401.690 1678.310 2402.870 ;
        RECT 1677.130 2223.290 1678.310 2224.470 ;
        RECT 1677.130 2221.690 1678.310 2222.870 ;
        RECT 1677.130 2043.290 1678.310 2044.470 ;
        RECT 1677.130 2041.690 1678.310 2042.870 ;
        RECT 1677.130 1863.290 1678.310 1864.470 ;
        RECT 1677.130 1861.690 1678.310 1862.870 ;
        RECT 1677.130 1683.290 1678.310 1684.470 ;
        RECT 1677.130 1681.690 1678.310 1682.870 ;
        RECT 1677.130 1503.290 1678.310 1504.470 ;
        RECT 1677.130 1501.690 1678.310 1502.870 ;
        RECT 1677.130 1323.290 1678.310 1324.470 ;
        RECT 1677.130 1321.690 1678.310 1322.870 ;
        RECT 1677.130 1143.290 1678.310 1144.470 ;
        RECT 1677.130 1141.690 1678.310 1142.870 ;
        RECT 1677.130 963.290 1678.310 964.470 ;
        RECT 1677.130 961.690 1678.310 962.870 ;
        RECT 1677.130 783.290 1678.310 784.470 ;
        RECT 1677.130 781.690 1678.310 782.870 ;
        RECT 1677.130 603.290 1678.310 604.470 ;
        RECT 1677.130 601.690 1678.310 602.870 ;
        RECT 1677.130 423.290 1678.310 424.470 ;
        RECT 1677.130 421.690 1678.310 422.870 ;
        RECT 1677.130 243.290 1678.310 244.470 ;
        RECT 1677.130 241.690 1678.310 242.870 ;
        RECT 1677.130 63.290 1678.310 64.470 ;
        RECT 1677.130 61.690 1678.310 62.870 ;
        RECT 1677.130 -30.510 1678.310 -29.330 ;
        RECT 1677.130 -32.110 1678.310 -30.930 ;
        RECT 1857.130 3550.610 1858.310 3551.790 ;
        RECT 1857.130 3549.010 1858.310 3550.190 ;
        RECT 1857.130 3483.290 1858.310 3484.470 ;
        RECT 1857.130 3481.690 1858.310 3482.870 ;
        RECT 1857.130 3303.290 1858.310 3304.470 ;
        RECT 1857.130 3301.690 1858.310 3302.870 ;
        RECT 1857.130 3123.290 1858.310 3124.470 ;
        RECT 1857.130 3121.690 1858.310 3122.870 ;
        RECT 1857.130 2943.290 1858.310 2944.470 ;
        RECT 1857.130 2941.690 1858.310 2942.870 ;
        RECT 1857.130 2763.290 1858.310 2764.470 ;
        RECT 1857.130 2761.690 1858.310 2762.870 ;
        RECT 1857.130 2583.290 1858.310 2584.470 ;
        RECT 1857.130 2581.690 1858.310 2582.870 ;
        RECT 1857.130 2403.290 1858.310 2404.470 ;
        RECT 1857.130 2401.690 1858.310 2402.870 ;
        RECT 1857.130 2223.290 1858.310 2224.470 ;
        RECT 1857.130 2221.690 1858.310 2222.870 ;
        RECT 1857.130 2043.290 1858.310 2044.470 ;
        RECT 1857.130 2041.690 1858.310 2042.870 ;
        RECT 1857.130 1863.290 1858.310 1864.470 ;
        RECT 1857.130 1861.690 1858.310 1862.870 ;
        RECT 1857.130 1683.290 1858.310 1684.470 ;
        RECT 1857.130 1681.690 1858.310 1682.870 ;
        RECT 1857.130 1503.290 1858.310 1504.470 ;
        RECT 1857.130 1501.690 1858.310 1502.870 ;
        RECT 1857.130 1323.290 1858.310 1324.470 ;
        RECT 1857.130 1321.690 1858.310 1322.870 ;
        RECT 1857.130 1143.290 1858.310 1144.470 ;
        RECT 1857.130 1141.690 1858.310 1142.870 ;
        RECT 1857.130 963.290 1858.310 964.470 ;
        RECT 1857.130 961.690 1858.310 962.870 ;
        RECT 1857.130 783.290 1858.310 784.470 ;
        RECT 1857.130 781.690 1858.310 782.870 ;
        RECT 1857.130 603.290 1858.310 604.470 ;
        RECT 1857.130 601.690 1858.310 602.870 ;
        RECT 1857.130 423.290 1858.310 424.470 ;
        RECT 1857.130 421.690 1858.310 422.870 ;
        RECT 1857.130 243.290 1858.310 244.470 ;
        RECT 1857.130 241.690 1858.310 242.870 ;
        RECT 1857.130 63.290 1858.310 64.470 ;
        RECT 1857.130 61.690 1858.310 62.870 ;
        RECT 1857.130 -30.510 1858.310 -29.330 ;
        RECT 1857.130 -32.110 1858.310 -30.930 ;
        RECT 2037.130 3550.610 2038.310 3551.790 ;
        RECT 2037.130 3549.010 2038.310 3550.190 ;
        RECT 2037.130 3483.290 2038.310 3484.470 ;
        RECT 2037.130 3481.690 2038.310 3482.870 ;
        RECT 2037.130 3303.290 2038.310 3304.470 ;
        RECT 2037.130 3301.690 2038.310 3302.870 ;
        RECT 2037.130 3123.290 2038.310 3124.470 ;
        RECT 2037.130 3121.690 2038.310 3122.870 ;
        RECT 2037.130 2943.290 2038.310 2944.470 ;
        RECT 2037.130 2941.690 2038.310 2942.870 ;
        RECT 2037.130 2763.290 2038.310 2764.470 ;
        RECT 2037.130 2761.690 2038.310 2762.870 ;
        RECT 2037.130 2583.290 2038.310 2584.470 ;
        RECT 2037.130 2581.690 2038.310 2582.870 ;
        RECT 2037.130 2403.290 2038.310 2404.470 ;
        RECT 2037.130 2401.690 2038.310 2402.870 ;
        RECT 2037.130 2223.290 2038.310 2224.470 ;
        RECT 2037.130 2221.690 2038.310 2222.870 ;
        RECT 2037.130 2043.290 2038.310 2044.470 ;
        RECT 2037.130 2041.690 2038.310 2042.870 ;
        RECT 2037.130 1863.290 2038.310 1864.470 ;
        RECT 2037.130 1861.690 2038.310 1862.870 ;
        RECT 2037.130 1683.290 2038.310 1684.470 ;
        RECT 2037.130 1681.690 2038.310 1682.870 ;
        RECT 2037.130 1503.290 2038.310 1504.470 ;
        RECT 2037.130 1501.690 2038.310 1502.870 ;
        RECT 2037.130 1323.290 2038.310 1324.470 ;
        RECT 2037.130 1321.690 2038.310 1322.870 ;
        RECT 2037.130 1143.290 2038.310 1144.470 ;
        RECT 2037.130 1141.690 2038.310 1142.870 ;
        RECT 2037.130 963.290 2038.310 964.470 ;
        RECT 2037.130 961.690 2038.310 962.870 ;
        RECT 2037.130 783.290 2038.310 784.470 ;
        RECT 2037.130 781.690 2038.310 782.870 ;
        RECT 2037.130 603.290 2038.310 604.470 ;
        RECT 2037.130 601.690 2038.310 602.870 ;
        RECT 2037.130 423.290 2038.310 424.470 ;
        RECT 2037.130 421.690 2038.310 422.870 ;
        RECT 2037.130 243.290 2038.310 244.470 ;
        RECT 2037.130 241.690 2038.310 242.870 ;
        RECT 2037.130 63.290 2038.310 64.470 ;
        RECT 2037.130 61.690 2038.310 62.870 ;
        RECT 2037.130 -30.510 2038.310 -29.330 ;
        RECT 2037.130 -32.110 2038.310 -30.930 ;
        RECT 2217.130 3550.610 2218.310 3551.790 ;
        RECT 2217.130 3549.010 2218.310 3550.190 ;
        RECT 2217.130 3483.290 2218.310 3484.470 ;
        RECT 2217.130 3481.690 2218.310 3482.870 ;
        RECT 2217.130 3303.290 2218.310 3304.470 ;
        RECT 2217.130 3301.690 2218.310 3302.870 ;
        RECT 2217.130 3123.290 2218.310 3124.470 ;
        RECT 2217.130 3121.690 2218.310 3122.870 ;
        RECT 2217.130 2943.290 2218.310 2944.470 ;
        RECT 2217.130 2941.690 2218.310 2942.870 ;
        RECT 2217.130 2763.290 2218.310 2764.470 ;
        RECT 2217.130 2761.690 2218.310 2762.870 ;
        RECT 2217.130 2583.290 2218.310 2584.470 ;
        RECT 2217.130 2581.690 2218.310 2582.870 ;
        RECT 2217.130 2403.290 2218.310 2404.470 ;
        RECT 2217.130 2401.690 2218.310 2402.870 ;
        RECT 2217.130 2223.290 2218.310 2224.470 ;
        RECT 2217.130 2221.690 2218.310 2222.870 ;
        RECT 2217.130 2043.290 2218.310 2044.470 ;
        RECT 2217.130 2041.690 2218.310 2042.870 ;
        RECT 2217.130 1863.290 2218.310 1864.470 ;
        RECT 2217.130 1861.690 2218.310 1862.870 ;
        RECT 2217.130 1683.290 2218.310 1684.470 ;
        RECT 2217.130 1681.690 2218.310 1682.870 ;
        RECT 2217.130 1503.290 2218.310 1504.470 ;
        RECT 2217.130 1501.690 2218.310 1502.870 ;
        RECT 2217.130 1323.290 2218.310 1324.470 ;
        RECT 2217.130 1321.690 2218.310 1322.870 ;
        RECT 2217.130 1143.290 2218.310 1144.470 ;
        RECT 2217.130 1141.690 2218.310 1142.870 ;
        RECT 2217.130 963.290 2218.310 964.470 ;
        RECT 2217.130 961.690 2218.310 962.870 ;
        RECT 2217.130 783.290 2218.310 784.470 ;
        RECT 2217.130 781.690 2218.310 782.870 ;
        RECT 2217.130 603.290 2218.310 604.470 ;
        RECT 2217.130 601.690 2218.310 602.870 ;
        RECT 2217.130 423.290 2218.310 424.470 ;
        RECT 2217.130 421.690 2218.310 422.870 ;
        RECT 2217.130 243.290 2218.310 244.470 ;
        RECT 2217.130 241.690 2218.310 242.870 ;
        RECT 2217.130 63.290 2218.310 64.470 ;
        RECT 2217.130 61.690 2218.310 62.870 ;
        RECT 2217.130 -30.510 2218.310 -29.330 ;
        RECT 2217.130 -32.110 2218.310 -30.930 ;
        RECT 2397.130 3550.610 2398.310 3551.790 ;
        RECT 2397.130 3549.010 2398.310 3550.190 ;
        RECT 2397.130 3483.290 2398.310 3484.470 ;
        RECT 2397.130 3481.690 2398.310 3482.870 ;
        RECT 2397.130 3303.290 2398.310 3304.470 ;
        RECT 2397.130 3301.690 2398.310 3302.870 ;
        RECT 2397.130 3123.290 2398.310 3124.470 ;
        RECT 2397.130 3121.690 2398.310 3122.870 ;
        RECT 2397.130 2943.290 2398.310 2944.470 ;
        RECT 2397.130 2941.690 2398.310 2942.870 ;
        RECT 2397.130 2763.290 2398.310 2764.470 ;
        RECT 2397.130 2761.690 2398.310 2762.870 ;
        RECT 2397.130 2583.290 2398.310 2584.470 ;
        RECT 2397.130 2581.690 2398.310 2582.870 ;
        RECT 2397.130 2403.290 2398.310 2404.470 ;
        RECT 2397.130 2401.690 2398.310 2402.870 ;
        RECT 2397.130 2223.290 2398.310 2224.470 ;
        RECT 2397.130 2221.690 2398.310 2222.870 ;
        RECT 2397.130 2043.290 2398.310 2044.470 ;
        RECT 2397.130 2041.690 2398.310 2042.870 ;
        RECT 2397.130 1863.290 2398.310 1864.470 ;
        RECT 2397.130 1861.690 2398.310 1862.870 ;
        RECT 2397.130 1683.290 2398.310 1684.470 ;
        RECT 2397.130 1681.690 2398.310 1682.870 ;
        RECT 2397.130 1503.290 2398.310 1504.470 ;
        RECT 2397.130 1501.690 2398.310 1502.870 ;
        RECT 2397.130 1323.290 2398.310 1324.470 ;
        RECT 2397.130 1321.690 2398.310 1322.870 ;
        RECT 2397.130 1143.290 2398.310 1144.470 ;
        RECT 2397.130 1141.690 2398.310 1142.870 ;
        RECT 2397.130 963.290 2398.310 964.470 ;
        RECT 2397.130 961.690 2398.310 962.870 ;
        RECT 2397.130 783.290 2398.310 784.470 ;
        RECT 2397.130 781.690 2398.310 782.870 ;
        RECT 2397.130 603.290 2398.310 604.470 ;
        RECT 2397.130 601.690 2398.310 602.870 ;
        RECT 2397.130 423.290 2398.310 424.470 ;
        RECT 2397.130 421.690 2398.310 422.870 ;
        RECT 2397.130 243.290 2398.310 244.470 ;
        RECT 2397.130 241.690 2398.310 242.870 ;
        RECT 2397.130 63.290 2398.310 64.470 ;
        RECT 2397.130 61.690 2398.310 62.870 ;
        RECT 2397.130 -30.510 2398.310 -29.330 ;
        RECT 2397.130 -32.110 2398.310 -30.930 ;
        RECT 2577.130 3550.610 2578.310 3551.790 ;
        RECT 2577.130 3549.010 2578.310 3550.190 ;
        RECT 2577.130 3483.290 2578.310 3484.470 ;
        RECT 2577.130 3481.690 2578.310 3482.870 ;
        RECT 2577.130 3303.290 2578.310 3304.470 ;
        RECT 2577.130 3301.690 2578.310 3302.870 ;
        RECT 2577.130 3123.290 2578.310 3124.470 ;
        RECT 2577.130 3121.690 2578.310 3122.870 ;
        RECT 2577.130 2943.290 2578.310 2944.470 ;
        RECT 2577.130 2941.690 2578.310 2942.870 ;
        RECT 2577.130 2763.290 2578.310 2764.470 ;
        RECT 2577.130 2761.690 2578.310 2762.870 ;
        RECT 2577.130 2583.290 2578.310 2584.470 ;
        RECT 2577.130 2581.690 2578.310 2582.870 ;
        RECT 2577.130 2403.290 2578.310 2404.470 ;
        RECT 2577.130 2401.690 2578.310 2402.870 ;
        RECT 2577.130 2223.290 2578.310 2224.470 ;
        RECT 2577.130 2221.690 2578.310 2222.870 ;
        RECT 2577.130 2043.290 2578.310 2044.470 ;
        RECT 2577.130 2041.690 2578.310 2042.870 ;
        RECT 2577.130 1863.290 2578.310 1864.470 ;
        RECT 2577.130 1861.690 2578.310 1862.870 ;
        RECT 2577.130 1683.290 2578.310 1684.470 ;
        RECT 2577.130 1681.690 2578.310 1682.870 ;
        RECT 2577.130 1503.290 2578.310 1504.470 ;
        RECT 2577.130 1501.690 2578.310 1502.870 ;
        RECT 2577.130 1323.290 2578.310 1324.470 ;
        RECT 2577.130 1321.690 2578.310 1322.870 ;
        RECT 2577.130 1143.290 2578.310 1144.470 ;
        RECT 2577.130 1141.690 2578.310 1142.870 ;
        RECT 2577.130 963.290 2578.310 964.470 ;
        RECT 2577.130 961.690 2578.310 962.870 ;
        RECT 2577.130 783.290 2578.310 784.470 ;
        RECT 2577.130 781.690 2578.310 782.870 ;
        RECT 2577.130 603.290 2578.310 604.470 ;
        RECT 2577.130 601.690 2578.310 602.870 ;
        RECT 2577.130 423.290 2578.310 424.470 ;
        RECT 2577.130 421.690 2578.310 422.870 ;
        RECT 2577.130 243.290 2578.310 244.470 ;
        RECT 2577.130 241.690 2578.310 242.870 ;
        RECT 2577.130 63.290 2578.310 64.470 ;
        RECT 2577.130 61.690 2578.310 62.870 ;
        RECT 2577.130 -30.510 2578.310 -29.330 ;
        RECT 2577.130 -32.110 2578.310 -30.930 ;
        RECT 2757.130 3550.610 2758.310 3551.790 ;
        RECT 2757.130 3549.010 2758.310 3550.190 ;
        RECT 2757.130 3483.290 2758.310 3484.470 ;
        RECT 2757.130 3481.690 2758.310 3482.870 ;
        RECT 2757.130 3303.290 2758.310 3304.470 ;
        RECT 2757.130 3301.690 2758.310 3302.870 ;
        RECT 2757.130 3123.290 2758.310 3124.470 ;
        RECT 2757.130 3121.690 2758.310 3122.870 ;
        RECT 2757.130 2943.290 2758.310 2944.470 ;
        RECT 2757.130 2941.690 2758.310 2942.870 ;
        RECT 2757.130 2763.290 2758.310 2764.470 ;
        RECT 2757.130 2761.690 2758.310 2762.870 ;
        RECT 2757.130 2583.290 2758.310 2584.470 ;
        RECT 2757.130 2581.690 2758.310 2582.870 ;
        RECT 2757.130 2403.290 2758.310 2404.470 ;
        RECT 2757.130 2401.690 2758.310 2402.870 ;
        RECT 2757.130 2223.290 2758.310 2224.470 ;
        RECT 2757.130 2221.690 2758.310 2222.870 ;
        RECT 2757.130 2043.290 2758.310 2044.470 ;
        RECT 2757.130 2041.690 2758.310 2042.870 ;
        RECT 2757.130 1863.290 2758.310 1864.470 ;
        RECT 2757.130 1861.690 2758.310 1862.870 ;
        RECT 2757.130 1683.290 2758.310 1684.470 ;
        RECT 2757.130 1681.690 2758.310 1682.870 ;
        RECT 2757.130 1503.290 2758.310 1504.470 ;
        RECT 2757.130 1501.690 2758.310 1502.870 ;
        RECT 2757.130 1323.290 2758.310 1324.470 ;
        RECT 2757.130 1321.690 2758.310 1322.870 ;
        RECT 2757.130 1143.290 2758.310 1144.470 ;
        RECT 2757.130 1141.690 2758.310 1142.870 ;
        RECT 2757.130 963.290 2758.310 964.470 ;
        RECT 2757.130 961.690 2758.310 962.870 ;
        RECT 2757.130 783.290 2758.310 784.470 ;
        RECT 2757.130 781.690 2758.310 782.870 ;
        RECT 2757.130 603.290 2758.310 604.470 ;
        RECT 2757.130 601.690 2758.310 602.870 ;
        RECT 2757.130 423.290 2758.310 424.470 ;
        RECT 2757.130 421.690 2758.310 422.870 ;
        RECT 2757.130 243.290 2758.310 244.470 ;
        RECT 2757.130 241.690 2758.310 242.870 ;
        RECT 2757.130 63.290 2758.310 64.470 ;
        RECT 2757.130 61.690 2758.310 62.870 ;
        RECT 2757.130 -30.510 2758.310 -29.330 ;
        RECT 2757.130 -32.110 2758.310 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3483.290 2956.290 3484.470 ;
        RECT 2955.110 3481.690 2956.290 3482.870 ;
        RECT 2955.110 3303.290 2956.290 3304.470 ;
        RECT 2955.110 3301.690 2956.290 3302.870 ;
        RECT 2955.110 3123.290 2956.290 3124.470 ;
        RECT 2955.110 3121.690 2956.290 3122.870 ;
        RECT 2955.110 2943.290 2956.290 2944.470 ;
        RECT 2955.110 2941.690 2956.290 2942.870 ;
        RECT 2955.110 2763.290 2956.290 2764.470 ;
        RECT 2955.110 2761.690 2956.290 2762.870 ;
        RECT 2955.110 2583.290 2956.290 2584.470 ;
        RECT 2955.110 2581.690 2956.290 2582.870 ;
        RECT 2955.110 2403.290 2956.290 2404.470 ;
        RECT 2955.110 2401.690 2956.290 2402.870 ;
        RECT 2955.110 2223.290 2956.290 2224.470 ;
        RECT 2955.110 2221.690 2956.290 2222.870 ;
        RECT 2955.110 2043.290 2956.290 2044.470 ;
        RECT 2955.110 2041.690 2956.290 2042.870 ;
        RECT 2955.110 1863.290 2956.290 1864.470 ;
        RECT 2955.110 1861.690 2956.290 1862.870 ;
        RECT 2955.110 1683.290 2956.290 1684.470 ;
        RECT 2955.110 1681.690 2956.290 1682.870 ;
        RECT 2955.110 1503.290 2956.290 1504.470 ;
        RECT 2955.110 1501.690 2956.290 1502.870 ;
        RECT 2955.110 1323.290 2956.290 1324.470 ;
        RECT 2955.110 1321.690 2956.290 1322.870 ;
        RECT 2955.110 1143.290 2956.290 1144.470 ;
        RECT 2955.110 1141.690 2956.290 1142.870 ;
        RECT 2955.110 963.290 2956.290 964.470 ;
        RECT 2955.110 961.690 2956.290 962.870 ;
        RECT 2955.110 783.290 2956.290 784.470 ;
        RECT 2955.110 781.690 2956.290 782.870 ;
        RECT 2955.110 603.290 2956.290 604.470 ;
        RECT 2955.110 601.690 2956.290 602.870 ;
        RECT 2955.110 423.290 2956.290 424.470 ;
        RECT 2955.110 421.690 2956.290 422.870 ;
        RECT 2955.110 243.290 2956.290 244.470 ;
        RECT 2955.110 241.690 2956.290 242.870 ;
        RECT 2955.110 63.290 2956.290 64.470 ;
        RECT 2955.110 61.690 2956.290 62.870 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.530 3551.850 -34.630 3551.910 ;
        RECT 56.270 3551.850 59.170 3551.910 ;
        RECT 236.270 3551.850 239.170 3551.910 ;
        RECT 416.270 3551.850 419.170 3551.910 ;
        RECT 596.270 3551.850 599.170 3551.910 ;
        RECT 776.270 3551.850 779.170 3551.910 ;
        RECT 956.270 3551.850 959.170 3551.910 ;
        RECT 1136.270 3551.850 1139.170 3551.910 ;
        RECT 1316.270 3551.850 1319.170 3551.910 ;
        RECT 1496.270 3551.850 1499.170 3551.910 ;
        RECT 1676.270 3551.850 1679.170 3551.910 ;
        RECT 1856.270 3551.850 1859.170 3551.910 ;
        RECT 2036.270 3551.850 2039.170 3551.910 ;
        RECT 2216.270 3551.850 2219.170 3551.910 ;
        RECT 2396.270 3551.850 2399.170 3551.910 ;
        RECT 2576.270 3551.850 2579.170 3551.910 ;
        RECT 2756.270 3551.850 2759.170 3551.910 ;
        RECT 2954.250 3551.850 2957.150 3551.910 ;
        RECT -37.530 3548.950 2957.150 3551.850 ;
        RECT -37.530 3548.890 -34.630 3548.950 ;
        RECT 56.270 3548.890 59.170 3548.950 ;
        RECT 236.270 3548.890 239.170 3548.950 ;
        RECT 416.270 3548.890 419.170 3548.950 ;
        RECT 596.270 3548.890 599.170 3548.950 ;
        RECT 776.270 3548.890 779.170 3548.950 ;
        RECT 956.270 3548.890 959.170 3548.950 ;
        RECT 1136.270 3548.890 1139.170 3548.950 ;
        RECT 1316.270 3548.890 1319.170 3548.950 ;
        RECT 1496.270 3548.890 1499.170 3548.950 ;
        RECT 1676.270 3548.890 1679.170 3548.950 ;
        RECT 1856.270 3548.890 1859.170 3548.950 ;
        RECT 2036.270 3548.890 2039.170 3548.950 ;
        RECT 2216.270 3548.890 2219.170 3548.950 ;
        RECT 2396.270 3548.890 2399.170 3548.950 ;
        RECT 2576.270 3548.890 2579.170 3548.950 ;
        RECT 2756.270 3548.890 2759.170 3548.950 ;
        RECT 2954.250 3548.890 2957.150 3548.950 ;
        RECT -37.530 3484.530 -34.630 3484.590 ;
        RECT 56.270 3484.530 59.170 3484.590 ;
        RECT 236.270 3484.530 239.170 3484.590 ;
        RECT 416.270 3484.530 419.170 3484.590 ;
        RECT 596.270 3484.530 599.170 3484.590 ;
        RECT 776.270 3484.530 779.170 3484.590 ;
        RECT 956.270 3484.530 959.170 3484.590 ;
        RECT 1136.270 3484.530 1139.170 3484.590 ;
        RECT 1316.270 3484.530 1319.170 3484.590 ;
        RECT 1496.270 3484.530 1499.170 3484.590 ;
        RECT 1676.270 3484.530 1679.170 3484.590 ;
        RECT 1856.270 3484.530 1859.170 3484.590 ;
        RECT 2036.270 3484.530 2039.170 3484.590 ;
        RECT 2216.270 3484.530 2219.170 3484.590 ;
        RECT 2396.270 3484.530 2399.170 3484.590 ;
        RECT 2576.270 3484.530 2579.170 3484.590 ;
        RECT 2756.270 3484.530 2759.170 3484.590 ;
        RECT 2954.250 3484.530 2957.150 3484.590 ;
        RECT -42.130 3481.630 2961.750 3484.530 ;
        RECT -37.530 3481.570 -34.630 3481.630 ;
        RECT 56.270 3481.570 59.170 3481.630 ;
        RECT 236.270 3481.570 239.170 3481.630 ;
        RECT 416.270 3481.570 419.170 3481.630 ;
        RECT 596.270 3481.570 599.170 3481.630 ;
        RECT 776.270 3481.570 779.170 3481.630 ;
        RECT 956.270 3481.570 959.170 3481.630 ;
        RECT 1136.270 3481.570 1139.170 3481.630 ;
        RECT 1316.270 3481.570 1319.170 3481.630 ;
        RECT 1496.270 3481.570 1499.170 3481.630 ;
        RECT 1676.270 3481.570 1679.170 3481.630 ;
        RECT 1856.270 3481.570 1859.170 3481.630 ;
        RECT 2036.270 3481.570 2039.170 3481.630 ;
        RECT 2216.270 3481.570 2219.170 3481.630 ;
        RECT 2396.270 3481.570 2399.170 3481.630 ;
        RECT 2576.270 3481.570 2579.170 3481.630 ;
        RECT 2756.270 3481.570 2759.170 3481.630 ;
        RECT 2954.250 3481.570 2957.150 3481.630 ;
        RECT -37.530 3304.530 -34.630 3304.590 ;
        RECT 56.270 3304.530 59.170 3304.590 ;
        RECT 236.270 3304.530 239.170 3304.590 ;
        RECT 416.270 3304.530 419.170 3304.590 ;
        RECT 596.270 3304.530 599.170 3304.590 ;
        RECT 776.270 3304.530 779.170 3304.590 ;
        RECT 956.270 3304.530 959.170 3304.590 ;
        RECT 1136.270 3304.530 1139.170 3304.590 ;
        RECT 1316.270 3304.530 1319.170 3304.590 ;
        RECT 1496.270 3304.530 1499.170 3304.590 ;
        RECT 1676.270 3304.530 1679.170 3304.590 ;
        RECT 1856.270 3304.530 1859.170 3304.590 ;
        RECT 2036.270 3304.530 2039.170 3304.590 ;
        RECT 2216.270 3304.530 2219.170 3304.590 ;
        RECT 2396.270 3304.530 2399.170 3304.590 ;
        RECT 2576.270 3304.530 2579.170 3304.590 ;
        RECT 2756.270 3304.530 2759.170 3304.590 ;
        RECT 2954.250 3304.530 2957.150 3304.590 ;
        RECT -42.130 3301.630 2961.750 3304.530 ;
        RECT -37.530 3301.570 -34.630 3301.630 ;
        RECT 56.270 3301.570 59.170 3301.630 ;
        RECT 236.270 3301.570 239.170 3301.630 ;
        RECT 416.270 3301.570 419.170 3301.630 ;
        RECT 596.270 3301.570 599.170 3301.630 ;
        RECT 776.270 3301.570 779.170 3301.630 ;
        RECT 956.270 3301.570 959.170 3301.630 ;
        RECT 1136.270 3301.570 1139.170 3301.630 ;
        RECT 1316.270 3301.570 1319.170 3301.630 ;
        RECT 1496.270 3301.570 1499.170 3301.630 ;
        RECT 1676.270 3301.570 1679.170 3301.630 ;
        RECT 1856.270 3301.570 1859.170 3301.630 ;
        RECT 2036.270 3301.570 2039.170 3301.630 ;
        RECT 2216.270 3301.570 2219.170 3301.630 ;
        RECT 2396.270 3301.570 2399.170 3301.630 ;
        RECT 2576.270 3301.570 2579.170 3301.630 ;
        RECT 2756.270 3301.570 2759.170 3301.630 ;
        RECT 2954.250 3301.570 2957.150 3301.630 ;
        RECT -37.530 3124.530 -34.630 3124.590 ;
        RECT 56.270 3124.530 59.170 3124.590 ;
        RECT 236.270 3124.530 239.170 3124.590 ;
        RECT 416.270 3124.530 419.170 3124.590 ;
        RECT 596.270 3124.530 599.170 3124.590 ;
        RECT 776.270 3124.530 779.170 3124.590 ;
        RECT 956.270 3124.530 959.170 3124.590 ;
        RECT 1136.270 3124.530 1139.170 3124.590 ;
        RECT 1316.270 3124.530 1319.170 3124.590 ;
        RECT 1496.270 3124.530 1499.170 3124.590 ;
        RECT 1676.270 3124.530 1679.170 3124.590 ;
        RECT 1856.270 3124.530 1859.170 3124.590 ;
        RECT 2036.270 3124.530 2039.170 3124.590 ;
        RECT 2216.270 3124.530 2219.170 3124.590 ;
        RECT 2396.270 3124.530 2399.170 3124.590 ;
        RECT 2576.270 3124.530 2579.170 3124.590 ;
        RECT 2756.270 3124.530 2759.170 3124.590 ;
        RECT 2954.250 3124.530 2957.150 3124.590 ;
        RECT -42.130 3121.630 2961.750 3124.530 ;
        RECT -37.530 3121.570 -34.630 3121.630 ;
        RECT 56.270 3121.570 59.170 3121.630 ;
        RECT 236.270 3121.570 239.170 3121.630 ;
        RECT 416.270 3121.570 419.170 3121.630 ;
        RECT 596.270 3121.570 599.170 3121.630 ;
        RECT 776.270 3121.570 779.170 3121.630 ;
        RECT 956.270 3121.570 959.170 3121.630 ;
        RECT 1136.270 3121.570 1139.170 3121.630 ;
        RECT 1316.270 3121.570 1319.170 3121.630 ;
        RECT 1496.270 3121.570 1499.170 3121.630 ;
        RECT 1676.270 3121.570 1679.170 3121.630 ;
        RECT 1856.270 3121.570 1859.170 3121.630 ;
        RECT 2036.270 3121.570 2039.170 3121.630 ;
        RECT 2216.270 3121.570 2219.170 3121.630 ;
        RECT 2396.270 3121.570 2399.170 3121.630 ;
        RECT 2576.270 3121.570 2579.170 3121.630 ;
        RECT 2756.270 3121.570 2759.170 3121.630 ;
        RECT 2954.250 3121.570 2957.150 3121.630 ;
        RECT -37.530 2944.530 -34.630 2944.590 ;
        RECT 56.270 2944.530 59.170 2944.590 ;
        RECT 236.270 2944.530 239.170 2944.590 ;
        RECT 416.270 2944.530 419.170 2944.590 ;
        RECT 596.270 2944.530 599.170 2944.590 ;
        RECT 776.270 2944.530 779.170 2944.590 ;
        RECT 956.270 2944.530 959.170 2944.590 ;
        RECT 1136.270 2944.530 1139.170 2944.590 ;
        RECT 1316.270 2944.530 1319.170 2944.590 ;
        RECT 1496.270 2944.530 1499.170 2944.590 ;
        RECT 1676.270 2944.530 1679.170 2944.590 ;
        RECT 1856.270 2944.530 1859.170 2944.590 ;
        RECT 2036.270 2944.530 2039.170 2944.590 ;
        RECT 2216.270 2944.530 2219.170 2944.590 ;
        RECT 2396.270 2944.530 2399.170 2944.590 ;
        RECT 2576.270 2944.530 2579.170 2944.590 ;
        RECT 2756.270 2944.530 2759.170 2944.590 ;
        RECT 2954.250 2944.530 2957.150 2944.590 ;
        RECT -42.130 2941.630 2961.750 2944.530 ;
        RECT -37.530 2941.570 -34.630 2941.630 ;
        RECT 56.270 2941.570 59.170 2941.630 ;
        RECT 236.270 2941.570 239.170 2941.630 ;
        RECT 416.270 2941.570 419.170 2941.630 ;
        RECT 596.270 2941.570 599.170 2941.630 ;
        RECT 776.270 2941.570 779.170 2941.630 ;
        RECT 956.270 2941.570 959.170 2941.630 ;
        RECT 1136.270 2941.570 1139.170 2941.630 ;
        RECT 1316.270 2941.570 1319.170 2941.630 ;
        RECT 1496.270 2941.570 1499.170 2941.630 ;
        RECT 1676.270 2941.570 1679.170 2941.630 ;
        RECT 1856.270 2941.570 1859.170 2941.630 ;
        RECT 2036.270 2941.570 2039.170 2941.630 ;
        RECT 2216.270 2941.570 2219.170 2941.630 ;
        RECT 2396.270 2941.570 2399.170 2941.630 ;
        RECT 2576.270 2941.570 2579.170 2941.630 ;
        RECT 2756.270 2941.570 2759.170 2941.630 ;
        RECT 2954.250 2941.570 2957.150 2941.630 ;
        RECT -37.530 2764.530 -34.630 2764.590 ;
        RECT 56.270 2764.530 59.170 2764.590 ;
        RECT 236.270 2764.530 239.170 2764.590 ;
        RECT 416.270 2764.530 419.170 2764.590 ;
        RECT 596.270 2764.530 599.170 2764.590 ;
        RECT 776.270 2764.530 779.170 2764.590 ;
        RECT 956.270 2764.530 959.170 2764.590 ;
        RECT 1136.270 2764.530 1139.170 2764.590 ;
        RECT 1316.270 2764.530 1319.170 2764.590 ;
        RECT 1496.270 2764.530 1499.170 2764.590 ;
        RECT 1676.270 2764.530 1679.170 2764.590 ;
        RECT 1856.270 2764.530 1859.170 2764.590 ;
        RECT 2036.270 2764.530 2039.170 2764.590 ;
        RECT 2216.270 2764.530 2219.170 2764.590 ;
        RECT 2396.270 2764.530 2399.170 2764.590 ;
        RECT 2576.270 2764.530 2579.170 2764.590 ;
        RECT 2756.270 2764.530 2759.170 2764.590 ;
        RECT 2954.250 2764.530 2957.150 2764.590 ;
        RECT -42.130 2761.630 2961.750 2764.530 ;
        RECT -37.530 2761.570 -34.630 2761.630 ;
        RECT 56.270 2761.570 59.170 2761.630 ;
        RECT 236.270 2761.570 239.170 2761.630 ;
        RECT 416.270 2761.570 419.170 2761.630 ;
        RECT 596.270 2761.570 599.170 2761.630 ;
        RECT 776.270 2761.570 779.170 2761.630 ;
        RECT 956.270 2761.570 959.170 2761.630 ;
        RECT 1136.270 2761.570 1139.170 2761.630 ;
        RECT 1316.270 2761.570 1319.170 2761.630 ;
        RECT 1496.270 2761.570 1499.170 2761.630 ;
        RECT 1676.270 2761.570 1679.170 2761.630 ;
        RECT 1856.270 2761.570 1859.170 2761.630 ;
        RECT 2036.270 2761.570 2039.170 2761.630 ;
        RECT 2216.270 2761.570 2219.170 2761.630 ;
        RECT 2396.270 2761.570 2399.170 2761.630 ;
        RECT 2576.270 2761.570 2579.170 2761.630 ;
        RECT 2756.270 2761.570 2759.170 2761.630 ;
        RECT 2954.250 2761.570 2957.150 2761.630 ;
        RECT -37.530 2584.530 -34.630 2584.590 ;
        RECT 56.270 2584.530 59.170 2584.590 ;
        RECT 236.270 2584.530 239.170 2584.590 ;
        RECT 416.270 2584.530 419.170 2584.590 ;
        RECT 596.270 2584.530 599.170 2584.590 ;
        RECT 776.270 2584.530 779.170 2584.590 ;
        RECT 956.270 2584.530 959.170 2584.590 ;
        RECT 1136.270 2584.530 1139.170 2584.590 ;
        RECT 1316.270 2584.530 1319.170 2584.590 ;
        RECT 1496.270 2584.530 1499.170 2584.590 ;
        RECT 1676.270 2584.530 1679.170 2584.590 ;
        RECT 1856.270 2584.530 1859.170 2584.590 ;
        RECT 2036.270 2584.530 2039.170 2584.590 ;
        RECT 2216.270 2584.530 2219.170 2584.590 ;
        RECT 2396.270 2584.530 2399.170 2584.590 ;
        RECT 2576.270 2584.530 2579.170 2584.590 ;
        RECT 2756.270 2584.530 2759.170 2584.590 ;
        RECT 2954.250 2584.530 2957.150 2584.590 ;
        RECT -42.130 2581.630 2961.750 2584.530 ;
        RECT -37.530 2581.570 -34.630 2581.630 ;
        RECT 56.270 2581.570 59.170 2581.630 ;
        RECT 236.270 2581.570 239.170 2581.630 ;
        RECT 416.270 2581.570 419.170 2581.630 ;
        RECT 596.270 2581.570 599.170 2581.630 ;
        RECT 776.270 2581.570 779.170 2581.630 ;
        RECT 956.270 2581.570 959.170 2581.630 ;
        RECT 1136.270 2581.570 1139.170 2581.630 ;
        RECT 1316.270 2581.570 1319.170 2581.630 ;
        RECT 1496.270 2581.570 1499.170 2581.630 ;
        RECT 1676.270 2581.570 1679.170 2581.630 ;
        RECT 1856.270 2581.570 1859.170 2581.630 ;
        RECT 2036.270 2581.570 2039.170 2581.630 ;
        RECT 2216.270 2581.570 2219.170 2581.630 ;
        RECT 2396.270 2581.570 2399.170 2581.630 ;
        RECT 2576.270 2581.570 2579.170 2581.630 ;
        RECT 2756.270 2581.570 2759.170 2581.630 ;
        RECT 2954.250 2581.570 2957.150 2581.630 ;
        RECT -37.530 2404.530 -34.630 2404.590 ;
        RECT 56.270 2404.530 59.170 2404.590 ;
        RECT 236.270 2404.530 239.170 2404.590 ;
        RECT 416.270 2404.530 419.170 2404.590 ;
        RECT 596.270 2404.530 599.170 2404.590 ;
        RECT 776.270 2404.530 779.170 2404.590 ;
        RECT 956.270 2404.530 959.170 2404.590 ;
        RECT 1136.270 2404.530 1139.170 2404.590 ;
        RECT 1316.270 2404.530 1319.170 2404.590 ;
        RECT 1496.270 2404.530 1499.170 2404.590 ;
        RECT 1676.270 2404.530 1679.170 2404.590 ;
        RECT 1856.270 2404.530 1859.170 2404.590 ;
        RECT 2036.270 2404.530 2039.170 2404.590 ;
        RECT 2216.270 2404.530 2219.170 2404.590 ;
        RECT 2396.270 2404.530 2399.170 2404.590 ;
        RECT 2576.270 2404.530 2579.170 2404.590 ;
        RECT 2756.270 2404.530 2759.170 2404.590 ;
        RECT 2954.250 2404.530 2957.150 2404.590 ;
        RECT -42.130 2401.630 2961.750 2404.530 ;
        RECT -37.530 2401.570 -34.630 2401.630 ;
        RECT 56.270 2401.570 59.170 2401.630 ;
        RECT 236.270 2401.570 239.170 2401.630 ;
        RECT 416.270 2401.570 419.170 2401.630 ;
        RECT 596.270 2401.570 599.170 2401.630 ;
        RECT 776.270 2401.570 779.170 2401.630 ;
        RECT 956.270 2401.570 959.170 2401.630 ;
        RECT 1136.270 2401.570 1139.170 2401.630 ;
        RECT 1316.270 2401.570 1319.170 2401.630 ;
        RECT 1496.270 2401.570 1499.170 2401.630 ;
        RECT 1676.270 2401.570 1679.170 2401.630 ;
        RECT 1856.270 2401.570 1859.170 2401.630 ;
        RECT 2036.270 2401.570 2039.170 2401.630 ;
        RECT 2216.270 2401.570 2219.170 2401.630 ;
        RECT 2396.270 2401.570 2399.170 2401.630 ;
        RECT 2576.270 2401.570 2579.170 2401.630 ;
        RECT 2756.270 2401.570 2759.170 2401.630 ;
        RECT 2954.250 2401.570 2957.150 2401.630 ;
        RECT -37.530 2224.530 -34.630 2224.590 ;
        RECT 56.270 2224.530 59.170 2224.590 ;
        RECT 236.270 2224.530 239.170 2224.590 ;
        RECT 416.270 2224.530 419.170 2224.590 ;
        RECT 596.270 2224.530 599.170 2224.590 ;
        RECT 776.270 2224.530 779.170 2224.590 ;
        RECT 956.270 2224.530 959.170 2224.590 ;
        RECT 1136.270 2224.530 1139.170 2224.590 ;
        RECT 1316.270 2224.530 1319.170 2224.590 ;
        RECT 1496.270 2224.530 1499.170 2224.590 ;
        RECT 1676.270 2224.530 1679.170 2224.590 ;
        RECT 1856.270 2224.530 1859.170 2224.590 ;
        RECT 2036.270 2224.530 2039.170 2224.590 ;
        RECT 2216.270 2224.530 2219.170 2224.590 ;
        RECT 2396.270 2224.530 2399.170 2224.590 ;
        RECT 2576.270 2224.530 2579.170 2224.590 ;
        RECT 2756.270 2224.530 2759.170 2224.590 ;
        RECT 2954.250 2224.530 2957.150 2224.590 ;
        RECT -42.130 2221.630 2961.750 2224.530 ;
        RECT -37.530 2221.570 -34.630 2221.630 ;
        RECT 56.270 2221.570 59.170 2221.630 ;
        RECT 236.270 2221.570 239.170 2221.630 ;
        RECT 416.270 2221.570 419.170 2221.630 ;
        RECT 596.270 2221.570 599.170 2221.630 ;
        RECT 776.270 2221.570 779.170 2221.630 ;
        RECT 956.270 2221.570 959.170 2221.630 ;
        RECT 1136.270 2221.570 1139.170 2221.630 ;
        RECT 1316.270 2221.570 1319.170 2221.630 ;
        RECT 1496.270 2221.570 1499.170 2221.630 ;
        RECT 1676.270 2221.570 1679.170 2221.630 ;
        RECT 1856.270 2221.570 1859.170 2221.630 ;
        RECT 2036.270 2221.570 2039.170 2221.630 ;
        RECT 2216.270 2221.570 2219.170 2221.630 ;
        RECT 2396.270 2221.570 2399.170 2221.630 ;
        RECT 2576.270 2221.570 2579.170 2221.630 ;
        RECT 2756.270 2221.570 2759.170 2221.630 ;
        RECT 2954.250 2221.570 2957.150 2221.630 ;
        RECT -37.530 2044.530 -34.630 2044.590 ;
        RECT 56.270 2044.530 59.170 2044.590 ;
        RECT 236.270 2044.530 239.170 2044.590 ;
        RECT 416.270 2044.530 419.170 2044.590 ;
        RECT 596.270 2044.530 599.170 2044.590 ;
        RECT 776.270 2044.530 779.170 2044.590 ;
        RECT 956.270 2044.530 959.170 2044.590 ;
        RECT 1136.270 2044.530 1139.170 2044.590 ;
        RECT 1316.270 2044.530 1319.170 2044.590 ;
        RECT 1496.270 2044.530 1499.170 2044.590 ;
        RECT 1676.270 2044.530 1679.170 2044.590 ;
        RECT 1856.270 2044.530 1859.170 2044.590 ;
        RECT 2036.270 2044.530 2039.170 2044.590 ;
        RECT 2216.270 2044.530 2219.170 2044.590 ;
        RECT 2396.270 2044.530 2399.170 2044.590 ;
        RECT 2576.270 2044.530 2579.170 2044.590 ;
        RECT 2756.270 2044.530 2759.170 2044.590 ;
        RECT 2954.250 2044.530 2957.150 2044.590 ;
        RECT -42.130 2041.630 2961.750 2044.530 ;
        RECT -37.530 2041.570 -34.630 2041.630 ;
        RECT 56.270 2041.570 59.170 2041.630 ;
        RECT 236.270 2041.570 239.170 2041.630 ;
        RECT 416.270 2041.570 419.170 2041.630 ;
        RECT 596.270 2041.570 599.170 2041.630 ;
        RECT 776.270 2041.570 779.170 2041.630 ;
        RECT 956.270 2041.570 959.170 2041.630 ;
        RECT 1136.270 2041.570 1139.170 2041.630 ;
        RECT 1316.270 2041.570 1319.170 2041.630 ;
        RECT 1496.270 2041.570 1499.170 2041.630 ;
        RECT 1676.270 2041.570 1679.170 2041.630 ;
        RECT 1856.270 2041.570 1859.170 2041.630 ;
        RECT 2036.270 2041.570 2039.170 2041.630 ;
        RECT 2216.270 2041.570 2219.170 2041.630 ;
        RECT 2396.270 2041.570 2399.170 2041.630 ;
        RECT 2576.270 2041.570 2579.170 2041.630 ;
        RECT 2756.270 2041.570 2759.170 2041.630 ;
        RECT 2954.250 2041.570 2957.150 2041.630 ;
        RECT -37.530 1864.530 -34.630 1864.590 ;
        RECT 56.270 1864.530 59.170 1864.590 ;
        RECT 236.270 1864.530 239.170 1864.590 ;
        RECT 416.270 1864.530 419.170 1864.590 ;
        RECT 596.270 1864.530 599.170 1864.590 ;
        RECT 776.270 1864.530 779.170 1864.590 ;
        RECT 956.270 1864.530 959.170 1864.590 ;
        RECT 1136.270 1864.530 1139.170 1864.590 ;
        RECT 1316.270 1864.530 1319.170 1864.590 ;
        RECT 1496.270 1864.530 1499.170 1864.590 ;
        RECT 1676.270 1864.530 1679.170 1864.590 ;
        RECT 1856.270 1864.530 1859.170 1864.590 ;
        RECT 2036.270 1864.530 2039.170 1864.590 ;
        RECT 2216.270 1864.530 2219.170 1864.590 ;
        RECT 2396.270 1864.530 2399.170 1864.590 ;
        RECT 2576.270 1864.530 2579.170 1864.590 ;
        RECT 2756.270 1864.530 2759.170 1864.590 ;
        RECT 2954.250 1864.530 2957.150 1864.590 ;
        RECT -42.130 1861.630 2961.750 1864.530 ;
        RECT -37.530 1861.570 -34.630 1861.630 ;
        RECT 56.270 1861.570 59.170 1861.630 ;
        RECT 236.270 1861.570 239.170 1861.630 ;
        RECT 416.270 1861.570 419.170 1861.630 ;
        RECT 596.270 1861.570 599.170 1861.630 ;
        RECT 776.270 1861.570 779.170 1861.630 ;
        RECT 956.270 1861.570 959.170 1861.630 ;
        RECT 1136.270 1861.570 1139.170 1861.630 ;
        RECT 1316.270 1861.570 1319.170 1861.630 ;
        RECT 1496.270 1861.570 1499.170 1861.630 ;
        RECT 1676.270 1861.570 1679.170 1861.630 ;
        RECT 1856.270 1861.570 1859.170 1861.630 ;
        RECT 2036.270 1861.570 2039.170 1861.630 ;
        RECT 2216.270 1861.570 2219.170 1861.630 ;
        RECT 2396.270 1861.570 2399.170 1861.630 ;
        RECT 2576.270 1861.570 2579.170 1861.630 ;
        RECT 2756.270 1861.570 2759.170 1861.630 ;
        RECT 2954.250 1861.570 2957.150 1861.630 ;
        RECT -37.530 1684.530 -34.630 1684.590 ;
        RECT 56.270 1684.530 59.170 1684.590 ;
        RECT 236.270 1684.530 239.170 1684.590 ;
        RECT 416.270 1684.530 419.170 1684.590 ;
        RECT 596.270 1684.530 599.170 1684.590 ;
        RECT 776.270 1684.530 779.170 1684.590 ;
        RECT 956.270 1684.530 959.170 1684.590 ;
        RECT 1136.270 1684.530 1139.170 1684.590 ;
        RECT 1316.270 1684.530 1319.170 1684.590 ;
        RECT 1496.270 1684.530 1499.170 1684.590 ;
        RECT 1676.270 1684.530 1679.170 1684.590 ;
        RECT 1856.270 1684.530 1859.170 1684.590 ;
        RECT 2036.270 1684.530 2039.170 1684.590 ;
        RECT 2216.270 1684.530 2219.170 1684.590 ;
        RECT 2396.270 1684.530 2399.170 1684.590 ;
        RECT 2576.270 1684.530 2579.170 1684.590 ;
        RECT 2756.270 1684.530 2759.170 1684.590 ;
        RECT 2954.250 1684.530 2957.150 1684.590 ;
        RECT -42.130 1681.630 2961.750 1684.530 ;
        RECT -37.530 1681.570 -34.630 1681.630 ;
        RECT 56.270 1681.570 59.170 1681.630 ;
        RECT 236.270 1681.570 239.170 1681.630 ;
        RECT 416.270 1681.570 419.170 1681.630 ;
        RECT 596.270 1681.570 599.170 1681.630 ;
        RECT 776.270 1681.570 779.170 1681.630 ;
        RECT 956.270 1681.570 959.170 1681.630 ;
        RECT 1136.270 1681.570 1139.170 1681.630 ;
        RECT 1316.270 1681.570 1319.170 1681.630 ;
        RECT 1496.270 1681.570 1499.170 1681.630 ;
        RECT 1676.270 1681.570 1679.170 1681.630 ;
        RECT 1856.270 1681.570 1859.170 1681.630 ;
        RECT 2036.270 1681.570 2039.170 1681.630 ;
        RECT 2216.270 1681.570 2219.170 1681.630 ;
        RECT 2396.270 1681.570 2399.170 1681.630 ;
        RECT 2576.270 1681.570 2579.170 1681.630 ;
        RECT 2756.270 1681.570 2759.170 1681.630 ;
        RECT 2954.250 1681.570 2957.150 1681.630 ;
        RECT -37.530 1504.530 -34.630 1504.590 ;
        RECT 56.270 1504.530 59.170 1504.590 ;
        RECT 236.270 1504.530 239.170 1504.590 ;
        RECT 416.270 1504.530 419.170 1504.590 ;
        RECT 596.270 1504.530 599.170 1504.590 ;
        RECT 776.270 1504.530 779.170 1504.590 ;
        RECT 956.270 1504.530 959.170 1504.590 ;
        RECT 1136.270 1504.530 1139.170 1504.590 ;
        RECT 1316.270 1504.530 1319.170 1504.590 ;
        RECT 1496.270 1504.530 1499.170 1504.590 ;
        RECT 1676.270 1504.530 1679.170 1504.590 ;
        RECT 1856.270 1504.530 1859.170 1504.590 ;
        RECT 2036.270 1504.530 2039.170 1504.590 ;
        RECT 2216.270 1504.530 2219.170 1504.590 ;
        RECT 2396.270 1504.530 2399.170 1504.590 ;
        RECT 2576.270 1504.530 2579.170 1504.590 ;
        RECT 2756.270 1504.530 2759.170 1504.590 ;
        RECT 2954.250 1504.530 2957.150 1504.590 ;
        RECT -42.130 1501.630 2961.750 1504.530 ;
        RECT -37.530 1501.570 -34.630 1501.630 ;
        RECT 56.270 1501.570 59.170 1501.630 ;
        RECT 236.270 1501.570 239.170 1501.630 ;
        RECT 416.270 1501.570 419.170 1501.630 ;
        RECT 596.270 1501.570 599.170 1501.630 ;
        RECT 776.270 1501.570 779.170 1501.630 ;
        RECT 956.270 1501.570 959.170 1501.630 ;
        RECT 1136.270 1501.570 1139.170 1501.630 ;
        RECT 1316.270 1501.570 1319.170 1501.630 ;
        RECT 1496.270 1501.570 1499.170 1501.630 ;
        RECT 1676.270 1501.570 1679.170 1501.630 ;
        RECT 1856.270 1501.570 1859.170 1501.630 ;
        RECT 2036.270 1501.570 2039.170 1501.630 ;
        RECT 2216.270 1501.570 2219.170 1501.630 ;
        RECT 2396.270 1501.570 2399.170 1501.630 ;
        RECT 2576.270 1501.570 2579.170 1501.630 ;
        RECT 2756.270 1501.570 2759.170 1501.630 ;
        RECT 2954.250 1501.570 2957.150 1501.630 ;
        RECT -37.530 1324.530 -34.630 1324.590 ;
        RECT 56.270 1324.530 59.170 1324.590 ;
        RECT 236.270 1324.530 239.170 1324.590 ;
        RECT 416.270 1324.530 419.170 1324.590 ;
        RECT 596.270 1324.530 599.170 1324.590 ;
        RECT 776.270 1324.530 779.170 1324.590 ;
        RECT 956.270 1324.530 959.170 1324.590 ;
        RECT 1136.270 1324.530 1139.170 1324.590 ;
        RECT 1316.270 1324.530 1319.170 1324.590 ;
        RECT 1496.270 1324.530 1499.170 1324.590 ;
        RECT 1676.270 1324.530 1679.170 1324.590 ;
        RECT 1856.270 1324.530 1859.170 1324.590 ;
        RECT 2036.270 1324.530 2039.170 1324.590 ;
        RECT 2216.270 1324.530 2219.170 1324.590 ;
        RECT 2396.270 1324.530 2399.170 1324.590 ;
        RECT 2576.270 1324.530 2579.170 1324.590 ;
        RECT 2756.270 1324.530 2759.170 1324.590 ;
        RECT 2954.250 1324.530 2957.150 1324.590 ;
        RECT -42.130 1321.630 2961.750 1324.530 ;
        RECT -37.530 1321.570 -34.630 1321.630 ;
        RECT 56.270 1321.570 59.170 1321.630 ;
        RECT 236.270 1321.570 239.170 1321.630 ;
        RECT 416.270 1321.570 419.170 1321.630 ;
        RECT 596.270 1321.570 599.170 1321.630 ;
        RECT 776.270 1321.570 779.170 1321.630 ;
        RECT 956.270 1321.570 959.170 1321.630 ;
        RECT 1136.270 1321.570 1139.170 1321.630 ;
        RECT 1316.270 1321.570 1319.170 1321.630 ;
        RECT 1496.270 1321.570 1499.170 1321.630 ;
        RECT 1676.270 1321.570 1679.170 1321.630 ;
        RECT 1856.270 1321.570 1859.170 1321.630 ;
        RECT 2036.270 1321.570 2039.170 1321.630 ;
        RECT 2216.270 1321.570 2219.170 1321.630 ;
        RECT 2396.270 1321.570 2399.170 1321.630 ;
        RECT 2576.270 1321.570 2579.170 1321.630 ;
        RECT 2756.270 1321.570 2759.170 1321.630 ;
        RECT 2954.250 1321.570 2957.150 1321.630 ;
        RECT -37.530 1144.530 -34.630 1144.590 ;
        RECT 56.270 1144.530 59.170 1144.590 ;
        RECT 236.270 1144.530 239.170 1144.590 ;
        RECT 416.270 1144.530 419.170 1144.590 ;
        RECT 596.270 1144.530 599.170 1144.590 ;
        RECT 776.270 1144.530 779.170 1144.590 ;
        RECT 956.270 1144.530 959.170 1144.590 ;
        RECT 1136.270 1144.530 1139.170 1144.590 ;
        RECT 1316.270 1144.530 1319.170 1144.590 ;
        RECT 1496.270 1144.530 1499.170 1144.590 ;
        RECT 1676.270 1144.530 1679.170 1144.590 ;
        RECT 1856.270 1144.530 1859.170 1144.590 ;
        RECT 2036.270 1144.530 2039.170 1144.590 ;
        RECT 2216.270 1144.530 2219.170 1144.590 ;
        RECT 2396.270 1144.530 2399.170 1144.590 ;
        RECT 2576.270 1144.530 2579.170 1144.590 ;
        RECT 2756.270 1144.530 2759.170 1144.590 ;
        RECT 2954.250 1144.530 2957.150 1144.590 ;
        RECT -42.130 1141.630 2961.750 1144.530 ;
        RECT -37.530 1141.570 -34.630 1141.630 ;
        RECT 56.270 1141.570 59.170 1141.630 ;
        RECT 236.270 1141.570 239.170 1141.630 ;
        RECT 416.270 1141.570 419.170 1141.630 ;
        RECT 596.270 1141.570 599.170 1141.630 ;
        RECT 776.270 1141.570 779.170 1141.630 ;
        RECT 956.270 1141.570 959.170 1141.630 ;
        RECT 1136.270 1141.570 1139.170 1141.630 ;
        RECT 1316.270 1141.570 1319.170 1141.630 ;
        RECT 1496.270 1141.570 1499.170 1141.630 ;
        RECT 1676.270 1141.570 1679.170 1141.630 ;
        RECT 1856.270 1141.570 1859.170 1141.630 ;
        RECT 2036.270 1141.570 2039.170 1141.630 ;
        RECT 2216.270 1141.570 2219.170 1141.630 ;
        RECT 2396.270 1141.570 2399.170 1141.630 ;
        RECT 2576.270 1141.570 2579.170 1141.630 ;
        RECT 2756.270 1141.570 2759.170 1141.630 ;
        RECT 2954.250 1141.570 2957.150 1141.630 ;
        RECT -37.530 964.530 -34.630 964.590 ;
        RECT 56.270 964.530 59.170 964.590 ;
        RECT 236.270 964.530 239.170 964.590 ;
        RECT 416.270 964.530 419.170 964.590 ;
        RECT 596.270 964.530 599.170 964.590 ;
        RECT 776.270 964.530 779.170 964.590 ;
        RECT 956.270 964.530 959.170 964.590 ;
        RECT 1136.270 964.530 1139.170 964.590 ;
        RECT 1316.270 964.530 1319.170 964.590 ;
        RECT 1496.270 964.530 1499.170 964.590 ;
        RECT 1676.270 964.530 1679.170 964.590 ;
        RECT 1856.270 964.530 1859.170 964.590 ;
        RECT 2036.270 964.530 2039.170 964.590 ;
        RECT 2216.270 964.530 2219.170 964.590 ;
        RECT 2396.270 964.530 2399.170 964.590 ;
        RECT 2576.270 964.530 2579.170 964.590 ;
        RECT 2756.270 964.530 2759.170 964.590 ;
        RECT 2954.250 964.530 2957.150 964.590 ;
        RECT -42.130 961.630 2961.750 964.530 ;
        RECT -37.530 961.570 -34.630 961.630 ;
        RECT 56.270 961.570 59.170 961.630 ;
        RECT 236.270 961.570 239.170 961.630 ;
        RECT 416.270 961.570 419.170 961.630 ;
        RECT 596.270 961.570 599.170 961.630 ;
        RECT 776.270 961.570 779.170 961.630 ;
        RECT 956.270 961.570 959.170 961.630 ;
        RECT 1136.270 961.570 1139.170 961.630 ;
        RECT 1316.270 961.570 1319.170 961.630 ;
        RECT 1496.270 961.570 1499.170 961.630 ;
        RECT 1676.270 961.570 1679.170 961.630 ;
        RECT 1856.270 961.570 1859.170 961.630 ;
        RECT 2036.270 961.570 2039.170 961.630 ;
        RECT 2216.270 961.570 2219.170 961.630 ;
        RECT 2396.270 961.570 2399.170 961.630 ;
        RECT 2576.270 961.570 2579.170 961.630 ;
        RECT 2756.270 961.570 2759.170 961.630 ;
        RECT 2954.250 961.570 2957.150 961.630 ;
        RECT -37.530 784.530 -34.630 784.590 ;
        RECT 56.270 784.530 59.170 784.590 ;
        RECT 236.270 784.530 239.170 784.590 ;
        RECT 416.270 784.530 419.170 784.590 ;
        RECT 596.270 784.530 599.170 784.590 ;
        RECT 776.270 784.530 779.170 784.590 ;
        RECT 956.270 784.530 959.170 784.590 ;
        RECT 1136.270 784.530 1139.170 784.590 ;
        RECT 1316.270 784.530 1319.170 784.590 ;
        RECT 1496.270 784.530 1499.170 784.590 ;
        RECT 1676.270 784.530 1679.170 784.590 ;
        RECT 1856.270 784.530 1859.170 784.590 ;
        RECT 2036.270 784.530 2039.170 784.590 ;
        RECT 2216.270 784.530 2219.170 784.590 ;
        RECT 2396.270 784.530 2399.170 784.590 ;
        RECT 2576.270 784.530 2579.170 784.590 ;
        RECT 2756.270 784.530 2759.170 784.590 ;
        RECT 2954.250 784.530 2957.150 784.590 ;
        RECT -42.130 781.630 2961.750 784.530 ;
        RECT -37.530 781.570 -34.630 781.630 ;
        RECT 56.270 781.570 59.170 781.630 ;
        RECT 236.270 781.570 239.170 781.630 ;
        RECT 416.270 781.570 419.170 781.630 ;
        RECT 596.270 781.570 599.170 781.630 ;
        RECT 776.270 781.570 779.170 781.630 ;
        RECT 956.270 781.570 959.170 781.630 ;
        RECT 1136.270 781.570 1139.170 781.630 ;
        RECT 1316.270 781.570 1319.170 781.630 ;
        RECT 1496.270 781.570 1499.170 781.630 ;
        RECT 1676.270 781.570 1679.170 781.630 ;
        RECT 1856.270 781.570 1859.170 781.630 ;
        RECT 2036.270 781.570 2039.170 781.630 ;
        RECT 2216.270 781.570 2219.170 781.630 ;
        RECT 2396.270 781.570 2399.170 781.630 ;
        RECT 2576.270 781.570 2579.170 781.630 ;
        RECT 2756.270 781.570 2759.170 781.630 ;
        RECT 2954.250 781.570 2957.150 781.630 ;
        RECT -37.530 604.530 -34.630 604.590 ;
        RECT 56.270 604.530 59.170 604.590 ;
        RECT 236.270 604.530 239.170 604.590 ;
        RECT 416.270 604.530 419.170 604.590 ;
        RECT 596.270 604.530 599.170 604.590 ;
        RECT 776.270 604.530 779.170 604.590 ;
        RECT 956.270 604.530 959.170 604.590 ;
        RECT 1136.270 604.530 1139.170 604.590 ;
        RECT 1316.270 604.530 1319.170 604.590 ;
        RECT 1496.270 604.530 1499.170 604.590 ;
        RECT 1676.270 604.530 1679.170 604.590 ;
        RECT 1856.270 604.530 1859.170 604.590 ;
        RECT 2036.270 604.530 2039.170 604.590 ;
        RECT 2216.270 604.530 2219.170 604.590 ;
        RECT 2396.270 604.530 2399.170 604.590 ;
        RECT 2576.270 604.530 2579.170 604.590 ;
        RECT 2756.270 604.530 2759.170 604.590 ;
        RECT 2954.250 604.530 2957.150 604.590 ;
        RECT -42.130 601.630 2961.750 604.530 ;
        RECT -37.530 601.570 -34.630 601.630 ;
        RECT 56.270 601.570 59.170 601.630 ;
        RECT 236.270 601.570 239.170 601.630 ;
        RECT 416.270 601.570 419.170 601.630 ;
        RECT 596.270 601.570 599.170 601.630 ;
        RECT 776.270 601.570 779.170 601.630 ;
        RECT 956.270 601.570 959.170 601.630 ;
        RECT 1136.270 601.570 1139.170 601.630 ;
        RECT 1316.270 601.570 1319.170 601.630 ;
        RECT 1496.270 601.570 1499.170 601.630 ;
        RECT 1676.270 601.570 1679.170 601.630 ;
        RECT 1856.270 601.570 1859.170 601.630 ;
        RECT 2036.270 601.570 2039.170 601.630 ;
        RECT 2216.270 601.570 2219.170 601.630 ;
        RECT 2396.270 601.570 2399.170 601.630 ;
        RECT 2576.270 601.570 2579.170 601.630 ;
        RECT 2756.270 601.570 2759.170 601.630 ;
        RECT 2954.250 601.570 2957.150 601.630 ;
        RECT -37.530 424.530 -34.630 424.590 ;
        RECT 56.270 424.530 59.170 424.590 ;
        RECT 236.270 424.530 239.170 424.590 ;
        RECT 416.270 424.530 419.170 424.590 ;
        RECT 596.270 424.530 599.170 424.590 ;
        RECT 776.270 424.530 779.170 424.590 ;
        RECT 956.270 424.530 959.170 424.590 ;
        RECT 1136.270 424.530 1139.170 424.590 ;
        RECT 1316.270 424.530 1319.170 424.590 ;
        RECT 1496.270 424.530 1499.170 424.590 ;
        RECT 1676.270 424.530 1679.170 424.590 ;
        RECT 1856.270 424.530 1859.170 424.590 ;
        RECT 2036.270 424.530 2039.170 424.590 ;
        RECT 2216.270 424.530 2219.170 424.590 ;
        RECT 2396.270 424.530 2399.170 424.590 ;
        RECT 2576.270 424.530 2579.170 424.590 ;
        RECT 2756.270 424.530 2759.170 424.590 ;
        RECT 2954.250 424.530 2957.150 424.590 ;
        RECT -42.130 421.630 2961.750 424.530 ;
        RECT -37.530 421.570 -34.630 421.630 ;
        RECT 56.270 421.570 59.170 421.630 ;
        RECT 236.270 421.570 239.170 421.630 ;
        RECT 416.270 421.570 419.170 421.630 ;
        RECT 596.270 421.570 599.170 421.630 ;
        RECT 776.270 421.570 779.170 421.630 ;
        RECT 956.270 421.570 959.170 421.630 ;
        RECT 1136.270 421.570 1139.170 421.630 ;
        RECT 1316.270 421.570 1319.170 421.630 ;
        RECT 1496.270 421.570 1499.170 421.630 ;
        RECT 1676.270 421.570 1679.170 421.630 ;
        RECT 1856.270 421.570 1859.170 421.630 ;
        RECT 2036.270 421.570 2039.170 421.630 ;
        RECT 2216.270 421.570 2219.170 421.630 ;
        RECT 2396.270 421.570 2399.170 421.630 ;
        RECT 2576.270 421.570 2579.170 421.630 ;
        RECT 2756.270 421.570 2759.170 421.630 ;
        RECT 2954.250 421.570 2957.150 421.630 ;
        RECT -37.530 244.530 -34.630 244.590 ;
        RECT 56.270 244.530 59.170 244.590 ;
        RECT 236.270 244.530 239.170 244.590 ;
        RECT 416.270 244.530 419.170 244.590 ;
        RECT 596.270 244.530 599.170 244.590 ;
        RECT 776.270 244.530 779.170 244.590 ;
        RECT 956.270 244.530 959.170 244.590 ;
        RECT 1136.270 244.530 1139.170 244.590 ;
        RECT 1316.270 244.530 1319.170 244.590 ;
        RECT 1496.270 244.530 1499.170 244.590 ;
        RECT 1676.270 244.530 1679.170 244.590 ;
        RECT 1856.270 244.530 1859.170 244.590 ;
        RECT 2036.270 244.530 2039.170 244.590 ;
        RECT 2216.270 244.530 2219.170 244.590 ;
        RECT 2396.270 244.530 2399.170 244.590 ;
        RECT 2576.270 244.530 2579.170 244.590 ;
        RECT 2756.270 244.530 2759.170 244.590 ;
        RECT 2954.250 244.530 2957.150 244.590 ;
        RECT -42.130 241.630 2961.750 244.530 ;
        RECT -37.530 241.570 -34.630 241.630 ;
        RECT 56.270 241.570 59.170 241.630 ;
        RECT 236.270 241.570 239.170 241.630 ;
        RECT 416.270 241.570 419.170 241.630 ;
        RECT 596.270 241.570 599.170 241.630 ;
        RECT 776.270 241.570 779.170 241.630 ;
        RECT 956.270 241.570 959.170 241.630 ;
        RECT 1136.270 241.570 1139.170 241.630 ;
        RECT 1316.270 241.570 1319.170 241.630 ;
        RECT 1496.270 241.570 1499.170 241.630 ;
        RECT 1676.270 241.570 1679.170 241.630 ;
        RECT 1856.270 241.570 1859.170 241.630 ;
        RECT 2036.270 241.570 2039.170 241.630 ;
        RECT 2216.270 241.570 2219.170 241.630 ;
        RECT 2396.270 241.570 2399.170 241.630 ;
        RECT 2576.270 241.570 2579.170 241.630 ;
        RECT 2756.270 241.570 2759.170 241.630 ;
        RECT 2954.250 241.570 2957.150 241.630 ;
        RECT -37.530 64.530 -34.630 64.590 ;
        RECT 56.270 64.530 59.170 64.590 ;
        RECT 236.270 64.530 239.170 64.590 ;
        RECT 416.270 64.530 419.170 64.590 ;
        RECT 596.270 64.530 599.170 64.590 ;
        RECT 776.270 64.530 779.170 64.590 ;
        RECT 956.270 64.530 959.170 64.590 ;
        RECT 1136.270 64.530 1139.170 64.590 ;
        RECT 1316.270 64.530 1319.170 64.590 ;
        RECT 1496.270 64.530 1499.170 64.590 ;
        RECT 1676.270 64.530 1679.170 64.590 ;
        RECT 1856.270 64.530 1859.170 64.590 ;
        RECT 2036.270 64.530 2039.170 64.590 ;
        RECT 2216.270 64.530 2219.170 64.590 ;
        RECT 2396.270 64.530 2399.170 64.590 ;
        RECT 2576.270 64.530 2579.170 64.590 ;
        RECT 2756.270 64.530 2759.170 64.590 ;
        RECT 2954.250 64.530 2957.150 64.590 ;
        RECT -42.130 61.630 2961.750 64.530 ;
        RECT -37.530 61.570 -34.630 61.630 ;
        RECT 56.270 61.570 59.170 61.630 ;
        RECT 236.270 61.570 239.170 61.630 ;
        RECT 416.270 61.570 419.170 61.630 ;
        RECT 596.270 61.570 599.170 61.630 ;
        RECT 776.270 61.570 779.170 61.630 ;
        RECT 956.270 61.570 959.170 61.630 ;
        RECT 1136.270 61.570 1139.170 61.630 ;
        RECT 1316.270 61.570 1319.170 61.630 ;
        RECT 1496.270 61.570 1499.170 61.630 ;
        RECT 1676.270 61.570 1679.170 61.630 ;
        RECT 1856.270 61.570 1859.170 61.630 ;
        RECT 2036.270 61.570 2039.170 61.630 ;
        RECT 2216.270 61.570 2219.170 61.630 ;
        RECT 2396.270 61.570 2399.170 61.630 ;
        RECT 2576.270 61.570 2579.170 61.630 ;
        RECT 2756.270 61.570 2759.170 61.630 ;
        RECT 2954.250 61.570 2957.150 61.630 ;
        RECT -37.530 -29.270 -34.630 -29.210 ;
        RECT 56.270 -29.270 59.170 -29.210 ;
        RECT 236.270 -29.270 239.170 -29.210 ;
        RECT 416.270 -29.270 419.170 -29.210 ;
        RECT 596.270 -29.270 599.170 -29.210 ;
        RECT 776.270 -29.270 779.170 -29.210 ;
        RECT 956.270 -29.270 959.170 -29.210 ;
        RECT 1136.270 -29.270 1139.170 -29.210 ;
        RECT 1316.270 -29.270 1319.170 -29.210 ;
        RECT 1496.270 -29.270 1499.170 -29.210 ;
        RECT 1676.270 -29.270 1679.170 -29.210 ;
        RECT 1856.270 -29.270 1859.170 -29.210 ;
        RECT 2036.270 -29.270 2039.170 -29.210 ;
        RECT 2216.270 -29.270 2219.170 -29.210 ;
        RECT 2396.270 -29.270 2399.170 -29.210 ;
        RECT 2576.270 -29.270 2579.170 -29.210 ;
        RECT 2756.270 -29.270 2759.170 -29.210 ;
        RECT 2954.250 -29.270 2957.150 -29.210 ;
        RECT -37.530 -32.170 2957.150 -29.270 ;
        RECT -37.530 -32.230 -34.630 -32.170 ;
        RECT 56.270 -32.230 59.170 -32.170 ;
        RECT 236.270 -32.230 239.170 -32.170 ;
        RECT 416.270 -32.230 419.170 -32.170 ;
        RECT 596.270 -32.230 599.170 -32.170 ;
        RECT 776.270 -32.230 779.170 -32.170 ;
        RECT 956.270 -32.230 959.170 -32.170 ;
        RECT 1136.270 -32.230 1139.170 -32.170 ;
        RECT 1316.270 -32.230 1319.170 -32.170 ;
        RECT 1496.270 -32.230 1499.170 -32.170 ;
        RECT 1676.270 -32.230 1679.170 -32.170 ;
        RECT 1856.270 -32.230 1859.170 -32.170 ;
        RECT 2036.270 -32.230 2039.170 -32.170 ;
        RECT 2216.270 -32.230 2219.170 -32.170 ;
        RECT 2396.270 -32.230 2399.170 -32.170 ;
        RECT 2576.270 -32.230 2579.170 -32.170 ;
        RECT 2756.270 -32.230 2759.170 -32.170 ;
        RECT 2954.250 -32.230 2957.150 -32.170 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.130 -36.770 -39.230 3556.450 ;
        RECT 146.270 -36.770 149.170 3556.450 ;
        RECT 326.270 -36.770 329.170 3556.450 ;
        RECT 506.270 -36.770 509.170 3556.450 ;
        RECT 686.270 -36.770 689.170 3556.450 ;
        RECT 866.270 -36.770 869.170 3556.450 ;
        RECT 1046.270 -36.770 1049.170 3556.450 ;
        RECT 1226.270 -36.770 1229.170 3556.450 ;
        RECT 1406.270 -36.770 1409.170 3556.450 ;
        RECT 1586.270 -36.770 1589.170 3556.450 ;
        RECT 1766.270 -36.770 1769.170 3556.450 ;
        RECT 1946.270 -36.770 1949.170 3556.450 ;
        RECT 2126.270 -36.770 2129.170 3556.450 ;
        RECT 2306.270 -36.770 2309.170 3556.450 ;
        RECT 2486.270 -36.770 2489.170 3556.450 ;
        RECT 2666.270 -36.770 2669.170 3556.450 ;
        RECT 2846.270 -36.770 2849.170 3556.450 ;
        RECT 2958.850 -36.770 2961.750 3556.450 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3393.290 -40.090 3394.470 ;
        RECT -41.270 3391.690 -40.090 3392.870 ;
        RECT -41.270 3213.290 -40.090 3214.470 ;
        RECT -41.270 3211.690 -40.090 3212.870 ;
        RECT -41.270 3033.290 -40.090 3034.470 ;
        RECT -41.270 3031.690 -40.090 3032.870 ;
        RECT -41.270 2853.290 -40.090 2854.470 ;
        RECT -41.270 2851.690 -40.090 2852.870 ;
        RECT -41.270 2673.290 -40.090 2674.470 ;
        RECT -41.270 2671.690 -40.090 2672.870 ;
        RECT -41.270 2493.290 -40.090 2494.470 ;
        RECT -41.270 2491.690 -40.090 2492.870 ;
        RECT -41.270 2313.290 -40.090 2314.470 ;
        RECT -41.270 2311.690 -40.090 2312.870 ;
        RECT -41.270 2133.290 -40.090 2134.470 ;
        RECT -41.270 2131.690 -40.090 2132.870 ;
        RECT -41.270 1953.290 -40.090 1954.470 ;
        RECT -41.270 1951.690 -40.090 1952.870 ;
        RECT -41.270 1773.290 -40.090 1774.470 ;
        RECT -41.270 1771.690 -40.090 1772.870 ;
        RECT -41.270 1593.290 -40.090 1594.470 ;
        RECT -41.270 1591.690 -40.090 1592.870 ;
        RECT -41.270 1413.290 -40.090 1414.470 ;
        RECT -41.270 1411.690 -40.090 1412.870 ;
        RECT -41.270 1233.290 -40.090 1234.470 ;
        RECT -41.270 1231.690 -40.090 1232.870 ;
        RECT -41.270 1053.290 -40.090 1054.470 ;
        RECT -41.270 1051.690 -40.090 1052.870 ;
        RECT -41.270 873.290 -40.090 874.470 ;
        RECT -41.270 871.690 -40.090 872.870 ;
        RECT -41.270 693.290 -40.090 694.470 ;
        RECT -41.270 691.690 -40.090 692.870 ;
        RECT -41.270 513.290 -40.090 514.470 ;
        RECT -41.270 511.690 -40.090 512.870 ;
        RECT -41.270 333.290 -40.090 334.470 ;
        RECT -41.270 331.690 -40.090 332.870 ;
        RECT -41.270 153.290 -40.090 154.470 ;
        RECT -41.270 151.690 -40.090 152.870 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 147.130 3555.210 148.310 3556.390 ;
        RECT 147.130 3553.610 148.310 3554.790 ;
        RECT 147.130 3393.290 148.310 3394.470 ;
        RECT 147.130 3391.690 148.310 3392.870 ;
        RECT 147.130 3213.290 148.310 3214.470 ;
        RECT 147.130 3211.690 148.310 3212.870 ;
        RECT 147.130 3033.290 148.310 3034.470 ;
        RECT 147.130 3031.690 148.310 3032.870 ;
        RECT 147.130 2853.290 148.310 2854.470 ;
        RECT 147.130 2851.690 148.310 2852.870 ;
        RECT 147.130 2673.290 148.310 2674.470 ;
        RECT 147.130 2671.690 148.310 2672.870 ;
        RECT 147.130 2493.290 148.310 2494.470 ;
        RECT 147.130 2491.690 148.310 2492.870 ;
        RECT 147.130 2313.290 148.310 2314.470 ;
        RECT 147.130 2311.690 148.310 2312.870 ;
        RECT 147.130 2133.290 148.310 2134.470 ;
        RECT 147.130 2131.690 148.310 2132.870 ;
        RECT 147.130 1953.290 148.310 1954.470 ;
        RECT 147.130 1951.690 148.310 1952.870 ;
        RECT 147.130 1773.290 148.310 1774.470 ;
        RECT 147.130 1771.690 148.310 1772.870 ;
        RECT 147.130 1593.290 148.310 1594.470 ;
        RECT 147.130 1591.690 148.310 1592.870 ;
        RECT 147.130 1413.290 148.310 1414.470 ;
        RECT 147.130 1411.690 148.310 1412.870 ;
        RECT 147.130 1233.290 148.310 1234.470 ;
        RECT 147.130 1231.690 148.310 1232.870 ;
        RECT 147.130 1053.290 148.310 1054.470 ;
        RECT 147.130 1051.690 148.310 1052.870 ;
        RECT 147.130 873.290 148.310 874.470 ;
        RECT 147.130 871.690 148.310 872.870 ;
        RECT 147.130 693.290 148.310 694.470 ;
        RECT 147.130 691.690 148.310 692.870 ;
        RECT 147.130 513.290 148.310 514.470 ;
        RECT 147.130 511.690 148.310 512.870 ;
        RECT 147.130 333.290 148.310 334.470 ;
        RECT 147.130 331.690 148.310 332.870 ;
        RECT 147.130 153.290 148.310 154.470 ;
        RECT 147.130 151.690 148.310 152.870 ;
        RECT 147.130 -35.110 148.310 -33.930 ;
        RECT 147.130 -36.710 148.310 -35.530 ;
        RECT 327.130 3555.210 328.310 3556.390 ;
        RECT 327.130 3553.610 328.310 3554.790 ;
        RECT 327.130 3393.290 328.310 3394.470 ;
        RECT 327.130 3391.690 328.310 3392.870 ;
        RECT 327.130 3213.290 328.310 3214.470 ;
        RECT 327.130 3211.690 328.310 3212.870 ;
        RECT 327.130 3033.290 328.310 3034.470 ;
        RECT 327.130 3031.690 328.310 3032.870 ;
        RECT 327.130 2853.290 328.310 2854.470 ;
        RECT 327.130 2851.690 328.310 2852.870 ;
        RECT 327.130 2673.290 328.310 2674.470 ;
        RECT 327.130 2671.690 328.310 2672.870 ;
        RECT 327.130 2493.290 328.310 2494.470 ;
        RECT 327.130 2491.690 328.310 2492.870 ;
        RECT 327.130 2313.290 328.310 2314.470 ;
        RECT 327.130 2311.690 328.310 2312.870 ;
        RECT 327.130 2133.290 328.310 2134.470 ;
        RECT 327.130 2131.690 328.310 2132.870 ;
        RECT 327.130 1953.290 328.310 1954.470 ;
        RECT 327.130 1951.690 328.310 1952.870 ;
        RECT 327.130 1773.290 328.310 1774.470 ;
        RECT 327.130 1771.690 328.310 1772.870 ;
        RECT 327.130 1593.290 328.310 1594.470 ;
        RECT 327.130 1591.690 328.310 1592.870 ;
        RECT 327.130 1413.290 328.310 1414.470 ;
        RECT 327.130 1411.690 328.310 1412.870 ;
        RECT 327.130 1233.290 328.310 1234.470 ;
        RECT 327.130 1231.690 328.310 1232.870 ;
        RECT 327.130 1053.290 328.310 1054.470 ;
        RECT 327.130 1051.690 328.310 1052.870 ;
        RECT 327.130 873.290 328.310 874.470 ;
        RECT 327.130 871.690 328.310 872.870 ;
        RECT 327.130 693.290 328.310 694.470 ;
        RECT 327.130 691.690 328.310 692.870 ;
        RECT 327.130 513.290 328.310 514.470 ;
        RECT 327.130 511.690 328.310 512.870 ;
        RECT 327.130 333.290 328.310 334.470 ;
        RECT 327.130 331.690 328.310 332.870 ;
        RECT 327.130 153.290 328.310 154.470 ;
        RECT 327.130 151.690 328.310 152.870 ;
        RECT 327.130 -35.110 328.310 -33.930 ;
        RECT 327.130 -36.710 328.310 -35.530 ;
        RECT 507.130 3555.210 508.310 3556.390 ;
        RECT 507.130 3553.610 508.310 3554.790 ;
        RECT 507.130 3393.290 508.310 3394.470 ;
        RECT 507.130 3391.690 508.310 3392.870 ;
        RECT 507.130 3213.290 508.310 3214.470 ;
        RECT 507.130 3211.690 508.310 3212.870 ;
        RECT 507.130 3033.290 508.310 3034.470 ;
        RECT 507.130 3031.690 508.310 3032.870 ;
        RECT 507.130 2853.290 508.310 2854.470 ;
        RECT 507.130 2851.690 508.310 2852.870 ;
        RECT 507.130 2673.290 508.310 2674.470 ;
        RECT 507.130 2671.690 508.310 2672.870 ;
        RECT 507.130 2493.290 508.310 2494.470 ;
        RECT 507.130 2491.690 508.310 2492.870 ;
        RECT 507.130 2313.290 508.310 2314.470 ;
        RECT 507.130 2311.690 508.310 2312.870 ;
        RECT 507.130 2133.290 508.310 2134.470 ;
        RECT 507.130 2131.690 508.310 2132.870 ;
        RECT 507.130 1953.290 508.310 1954.470 ;
        RECT 507.130 1951.690 508.310 1952.870 ;
        RECT 507.130 1773.290 508.310 1774.470 ;
        RECT 507.130 1771.690 508.310 1772.870 ;
        RECT 507.130 1593.290 508.310 1594.470 ;
        RECT 507.130 1591.690 508.310 1592.870 ;
        RECT 507.130 1413.290 508.310 1414.470 ;
        RECT 507.130 1411.690 508.310 1412.870 ;
        RECT 507.130 1233.290 508.310 1234.470 ;
        RECT 507.130 1231.690 508.310 1232.870 ;
        RECT 507.130 1053.290 508.310 1054.470 ;
        RECT 507.130 1051.690 508.310 1052.870 ;
        RECT 507.130 873.290 508.310 874.470 ;
        RECT 507.130 871.690 508.310 872.870 ;
        RECT 507.130 693.290 508.310 694.470 ;
        RECT 507.130 691.690 508.310 692.870 ;
        RECT 507.130 513.290 508.310 514.470 ;
        RECT 507.130 511.690 508.310 512.870 ;
        RECT 507.130 333.290 508.310 334.470 ;
        RECT 507.130 331.690 508.310 332.870 ;
        RECT 507.130 153.290 508.310 154.470 ;
        RECT 507.130 151.690 508.310 152.870 ;
        RECT 507.130 -35.110 508.310 -33.930 ;
        RECT 507.130 -36.710 508.310 -35.530 ;
        RECT 687.130 3555.210 688.310 3556.390 ;
        RECT 687.130 3553.610 688.310 3554.790 ;
        RECT 687.130 3393.290 688.310 3394.470 ;
        RECT 687.130 3391.690 688.310 3392.870 ;
        RECT 687.130 3213.290 688.310 3214.470 ;
        RECT 687.130 3211.690 688.310 3212.870 ;
        RECT 687.130 3033.290 688.310 3034.470 ;
        RECT 687.130 3031.690 688.310 3032.870 ;
        RECT 687.130 2853.290 688.310 2854.470 ;
        RECT 687.130 2851.690 688.310 2852.870 ;
        RECT 687.130 2673.290 688.310 2674.470 ;
        RECT 687.130 2671.690 688.310 2672.870 ;
        RECT 687.130 2493.290 688.310 2494.470 ;
        RECT 687.130 2491.690 688.310 2492.870 ;
        RECT 687.130 2313.290 688.310 2314.470 ;
        RECT 687.130 2311.690 688.310 2312.870 ;
        RECT 687.130 2133.290 688.310 2134.470 ;
        RECT 687.130 2131.690 688.310 2132.870 ;
        RECT 687.130 1953.290 688.310 1954.470 ;
        RECT 687.130 1951.690 688.310 1952.870 ;
        RECT 687.130 1773.290 688.310 1774.470 ;
        RECT 687.130 1771.690 688.310 1772.870 ;
        RECT 687.130 1593.290 688.310 1594.470 ;
        RECT 687.130 1591.690 688.310 1592.870 ;
        RECT 687.130 1413.290 688.310 1414.470 ;
        RECT 687.130 1411.690 688.310 1412.870 ;
        RECT 687.130 1233.290 688.310 1234.470 ;
        RECT 687.130 1231.690 688.310 1232.870 ;
        RECT 687.130 1053.290 688.310 1054.470 ;
        RECT 687.130 1051.690 688.310 1052.870 ;
        RECT 687.130 873.290 688.310 874.470 ;
        RECT 687.130 871.690 688.310 872.870 ;
        RECT 687.130 693.290 688.310 694.470 ;
        RECT 687.130 691.690 688.310 692.870 ;
        RECT 687.130 513.290 688.310 514.470 ;
        RECT 687.130 511.690 688.310 512.870 ;
        RECT 687.130 333.290 688.310 334.470 ;
        RECT 687.130 331.690 688.310 332.870 ;
        RECT 687.130 153.290 688.310 154.470 ;
        RECT 687.130 151.690 688.310 152.870 ;
        RECT 687.130 -35.110 688.310 -33.930 ;
        RECT 687.130 -36.710 688.310 -35.530 ;
        RECT 867.130 3555.210 868.310 3556.390 ;
        RECT 867.130 3553.610 868.310 3554.790 ;
        RECT 867.130 3393.290 868.310 3394.470 ;
        RECT 867.130 3391.690 868.310 3392.870 ;
        RECT 867.130 3213.290 868.310 3214.470 ;
        RECT 867.130 3211.690 868.310 3212.870 ;
        RECT 867.130 3033.290 868.310 3034.470 ;
        RECT 867.130 3031.690 868.310 3032.870 ;
        RECT 867.130 2853.290 868.310 2854.470 ;
        RECT 867.130 2851.690 868.310 2852.870 ;
        RECT 867.130 2673.290 868.310 2674.470 ;
        RECT 867.130 2671.690 868.310 2672.870 ;
        RECT 867.130 2493.290 868.310 2494.470 ;
        RECT 867.130 2491.690 868.310 2492.870 ;
        RECT 867.130 2313.290 868.310 2314.470 ;
        RECT 867.130 2311.690 868.310 2312.870 ;
        RECT 867.130 2133.290 868.310 2134.470 ;
        RECT 867.130 2131.690 868.310 2132.870 ;
        RECT 867.130 1953.290 868.310 1954.470 ;
        RECT 867.130 1951.690 868.310 1952.870 ;
        RECT 867.130 1773.290 868.310 1774.470 ;
        RECT 867.130 1771.690 868.310 1772.870 ;
        RECT 867.130 1593.290 868.310 1594.470 ;
        RECT 867.130 1591.690 868.310 1592.870 ;
        RECT 867.130 1413.290 868.310 1414.470 ;
        RECT 867.130 1411.690 868.310 1412.870 ;
        RECT 867.130 1233.290 868.310 1234.470 ;
        RECT 867.130 1231.690 868.310 1232.870 ;
        RECT 867.130 1053.290 868.310 1054.470 ;
        RECT 867.130 1051.690 868.310 1052.870 ;
        RECT 867.130 873.290 868.310 874.470 ;
        RECT 867.130 871.690 868.310 872.870 ;
        RECT 867.130 693.290 868.310 694.470 ;
        RECT 867.130 691.690 868.310 692.870 ;
        RECT 867.130 513.290 868.310 514.470 ;
        RECT 867.130 511.690 868.310 512.870 ;
        RECT 867.130 333.290 868.310 334.470 ;
        RECT 867.130 331.690 868.310 332.870 ;
        RECT 867.130 153.290 868.310 154.470 ;
        RECT 867.130 151.690 868.310 152.870 ;
        RECT 867.130 -35.110 868.310 -33.930 ;
        RECT 867.130 -36.710 868.310 -35.530 ;
        RECT 1047.130 3555.210 1048.310 3556.390 ;
        RECT 1047.130 3553.610 1048.310 3554.790 ;
        RECT 1047.130 3393.290 1048.310 3394.470 ;
        RECT 1047.130 3391.690 1048.310 3392.870 ;
        RECT 1047.130 3213.290 1048.310 3214.470 ;
        RECT 1047.130 3211.690 1048.310 3212.870 ;
        RECT 1047.130 3033.290 1048.310 3034.470 ;
        RECT 1047.130 3031.690 1048.310 3032.870 ;
        RECT 1047.130 2853.290 1048.310 2854.470 ;
        RECT 1047.130 2851.690 1048.310 2852.870 ;
        RECT 1047.130 2673.290 1048.310 2674.470 ;
        RECT 1047.130 2671.690 1048.310 2672.870 ;
        RECT 1047.130 2493.290 1048.310 2494.470 ;
        RECT 1047.130 2491.690 1048.310 2492.870 ;
        RECT 1047.130 2313.290 1048.310 2314.470 ;
        RECT 1047.130 2311.690 1048.310 2312.870 ;
        RECT 1047.130 2133.290 1048.310 2134.470 ;
        RECT 1047.130 2131.690 1048.310 2132.870 ;
        RECT 1047.130 1953.290 1048.310 1954.470 ;
        RECT 1047.130 1951.690 1048.310 1952.870 ;
        RECT 1047.130 1773.290 1048.310 1774.470 ;
        RECT 1047.130 1771.690 1048.310 1772.870 ;
        RECT 1047.130 1593.290 1048.310 1594.470 ;
        RECT 1047.130 1591.690 1048.310 1592.870 ;
        RECT 1047.130 1413.290 1048.310 1414.470 ;
        RECT 1047.130 1411.690 1048.310 1412.870 ;
        RECT 1047.130 1233.290 1048.310 1234.470 ;
        RECT 1047.130 1231.690 1048.310 1232.870 ;
        RECT 1047.130 1053.290 1048.310 1054.470 ;
        RECT 1047.130 1051.690 1048.310 1052.870 ;
        RECT 1047.130 873.290 1048.310 874.470 ;
        RECT 1047.130 871.690 1048.310 872.870 ;
        RECT 1047.130 693.290 1048.310 694.470 ;
        RECT 1047.130 691.690 1048.310 692.870 ;
        RECT 1047.130 513.290 1048.310 514.470 ;
        RECT 1047.130 511.690 1048.310 512.870 ;
        RECT 1047.130 333.290 1048.310 334.470 ;
        RECT 1047.130 331.690 1048.310 332.870 ;
        RECT 1047.130 153.290 1048.310 154.470 ;
        RECT 1047.130 151.690 1048.310 152.870 ;
        RECT 1047.130 -35.110 1048.310 -33.930 ;
        RECT 1047.130 -36.710 1048.310 -35.530 ;
        RECT 1227.130 3555.210 1228.310 3556.390 ;
        RECT 1227.130 3553.610 1228.310 3554.790 ;
        RECT 1227.130 3393.290 1228.310 3394.470 ;
        RECT 1227.130 3391.690 1228.310 3392.870 ;
        RECT 1227.130 3213.290 1228.310 3214.470 ;
        RECT 1227.130 3211.690 1228.310 3212.870 ;
        RECT 1227.130 3033.290 1228.310 3034.470 ;
        RECT 1227.130 3031.690 1228.310 3032.870 ;
        RECT 1227.130 2853.290 1228.310 2854.470 ;
        RECT 1227.130 2851.690 1228.310 2852.870 ;
        RECT 1227.130 2673.290 1228.310 2674.470 ;
        RECT 1227.130 2671.690 1228.310 2672.870 ;
        RECT 1227.130 2493.290 1228.310 2494.470 ;
        RECT 1227.130 2491.690 1228.310 2492.870 ;
        RECT 1227.130 2313.290 1228.310 2314.470 ;
        RECT 1227.130 2311.690 1228.310 2312.870 ;
        RECT 1227.130 2133.290 1228.310 2134.470 ;
        RECT 1227.130 2131.690 1228.310 2132.870 ;
        RECT 1227.130 1953.290 1228.310 1954.470 ;
        RECT 1227.130 1951.690 1228.310 1952.870 ;
        RECT 1227.130 1773.290 1228.310 1774.470 ;
        RECT 1227.130 1771.690 1228.310 1772.870 ;
        RECT 1227.130 1593.290 1228.310 1594.470 ;
        RECT 1227.130 1591.690 1228.310 1592.870 ;
        RECT 1227.130 1413.290 1228.310 1414.470 ;
        RECT 1227.130 1411.690 1228.310 1412.870 ;
        RECT 1227.130 1233.290 1228.310 1234.470 ;
        RECT 1227.130 1231.690 1228.310 1232.870 ;
        RECT 1227.130 1053.290 1228.310 1054.470 ;
        RECT 1227.130 1051.690 1228.310 1052.870 ;
        RECT 1227.130 873.290 1228.310 874.470 ;
        RECT 1227.130 871.690 1228.310 872.870 ;
        RECT 1227.130 693.290 1228.310 694.470 ;
        RECT 1227.130 691.690 1228.310 692.870 ;
        RECT 1227.130 513.290 1228.310 514.470 ;
        RECT 1227.130 511.690 1228.310 512.870 ;
        RECT 1227.130 333.290 1228.310 334.470 ;
        RECT 1227.130 331.690 1228.310 332.870 ;
        RECT 1227.130 153.290 1228.310 154.470 ;
        RECT 1227.130 151.690 1228.310 152.870 ;
        RECT 1227.130 -35.110 1228.310 -33.930 ;
        RECT 1227.130 -36.710 1228.310 -35.530 ;
        RECT 1407.130 3555.210 1408.310 3556.390 ;
        RECT 1407.130 3553.610 1408.310 3554.790 ;
        RECT 1407.130 3393.290 1408.310 3394.470 ;
        RECT 1407.130 3391.690 1408.310 3392.870 ;
        RECT 1407.130 3213.290 1408.310 3214.470 ;
        RECT 1407.130 3211.690 1408.310 3212.870 ;
        RECT 1407.130 3033.290 1408.310 3034.470 ;
        RECT 1407.130 3031.690 1408.310 3032.870 ;
        RECT 1407.130 2853.290 1408.310 2854.470 ;
        RECT 1407.130 2851.690 1408.310 2852.870 ;
        RECT 1407.130 2673.290 1408.310 2674.470 ;
        RECT 1407.130 2671.690 1408.310 2672.870 ;
        RECT 1407.130 2493.290 1408.310 2494.470 ;
        RECT 1407.130 2491.690 1408.310 2492.870 ;
        RECT 1407.130 2313.290 1408.310 2314.470 ;
        RECT 1407.130 2311.690 1408.310 2312.870 ;
        RECT 1407.130 2133.290 1408.310 2134.470 ;
        RECT 1407.130 2131.690 1408.310 2132.870 ;
        RECT 1407.130 1953.290 1408.310 1954.470 ;
        RECT 1407.130 1951.690 1408.310 1952.870 ;
        RECT 1407.130 1773.290 1408.310 1774.470 ;
        RECT 1407.130 1771.690 1408.310 1772.870 ;
        RECT 1407.130 1593.290 1408.310 1594.470 ;
        RECT 1407.130 1591.690 1408.310 1592.870 ;
        RECT 1407.130 1413.290 1408.310 1414.470 ;
        RECT 1407.130 1411.690 1408.310 1412.870 ;
        RECT 1407.130 1233.290 1408.310 1234.470 ;
        RECT 1407.130 1231.690 1408.310 1232.870 ;
        RECT 1407.130 1053.290 1408.310 1054.470 ;
        RECT 1407.130 1051.690 1408.310 1052.870 ;
        RECT 1407.130 873.290 1408.310 874.470 ;
        RECT 1407.130 871.690 1408.310 872.870 ;
        RECT 1407.130 693.290 1408.310 694.470 ;
        RECT 1407.130 691.690 1408.310 692.870 ;
        RECT 1407.130 513.290 1408.310 514.470 ;
        RECT 1407.130 511.690 1408.310 512.870 ;
        RECT 1407.130 333.290 1408.310 334.470 ;
        RECT 1407.130 331.690 1408.310 332.870 ;
        RECT 1407.130 153.290 1408.310 154.470 ;
        RECT 1407.130 151.690 1408.310 152.870 ;
        RECT 1407.130 -35.110 1408.310 -33.930 ;
        RECT 1407.130 -36.710 1408.310 -35.530 ;
        RECT 1587.130 3555.210 1588.310 3556.390 ;
        RECT 1587.130 3553.610 1588.310 3554.790 ;
        RECT 1587.130 3393.290 1588.310 3394.470 ;
        RECT 1587.130 3391.690 1588.310 3392.870 ;
        RECT 1587.130 3213.290 1588.310 3214.470 ;
        RECT 1587.130 3211.690 1588.310 3212.870 ;
        RECT 1587.130 3033.290 1588.310 3034.470 ;
        RECT 1587.130 3031.690 1588.310 3032.870 ;
        RECT 1587.130 2853.290 1588.310 2854.470 ;
        RECT 1587.130 2851.690 1588.310 2852.870 ;
        RECT 1587.130 2673.290 1588.310 2674.470 ;
        RECT 1587.130 2671.690 1588.310 2672.870 ;
        RECT 1587.130 2493.290 1588.310 2494.470 ;
        RECT 1587.130 2491.690 1588.310 2492.870 ;
        RECT 1587.130 2313.290 1588.310 2314.470 ;
        RECT 1587.130 2311.690 1588.310 2312.870 ;
        RECT 1587.130 2133.290 1588.310 2134.470 ;
        RECT 1587.130 2131.690 1588.310 2132.870 ;
        RECT 1587.130 1953.290 1588.310 1954.470 ;
        RECT 1587.130 1951.690 1588.310 1952.870 ;
        RECT 1587.130 1773.290 1588.310 1774.470 ;
        RECT 1587.130 1771.690 1588.310 1772.870 ;
        RECT 1587.130 1593.290 1588.310 1594.470 ;
        RECT 1587.130 1591.690 1588.310 1592.870 ;
        RECT 1587.130 1413.290 1588.310 1414.470 ;
        RECT 1587.130 1411.690 1588.310 1412.870 ;
        RECT 1587.130 1233.290 1588.310 1234.470 ;
        RECT 1587.130 1231.690 1588.310 1232.870 ;
        RECT 1587.130 1053.290 1588.310 1054.470 ;
        RECT 1587.130 1051.690 1588.310 1052.870 ;
        RECT 1587.130 873.290 1588.310 874.470 ;
        RECT 1587.130 871.690 1588.310 872.870 ;
        RECT 1587.130 693.290 1588.310 694.470 ;
        RECT 1587.130 691.690 1588.310 692.870 ;
        RECT 1587.130 513.290 1588.310 514.470 ;
        RECT 1587.130 511.690 1588.310 512.870 ;
        RECT 1587.130 333.290 1588.310 334.470 ;
        RECT 1587.130 331.690 1588.310 332.870 ;
        RECT 1587.130 153.290 1588.310 154.470 ;
        RECT 1587.130 151.690 1588.310 152.870 ;
        RECT 1587.130 -35.110 1588.310 -33.930 ;
        RECT 1587.130 -36.710 1588.310 -35.530 ;
        RECT 1767.130 3555.210 1768.310 3556.390 ;
        RECT 1767.130 3553.610 1768.310 3554.790 ;
        RECT 1767.130 3393.290 1768.310 3394.470 ;
        RECT 1767.130 3391.690 1768.310 3392.870 ;
        RECT 1767.130 3213.290 1768.310 3214.470 ;
        RECT 1767.130 3211.690 1768.310 3212.870 ;
        RECT 1767.130 3033.290 1768.310 3034.470 ;
        RECT 1767.130 3031.690 1768.310 3032.870 ;
        RECT 1767.130 2853.290 1768.310 2854.470 ;
        RECT 1767.130 2851.690 1768.310 2852.870 ;
        RECT 1767.130 2673.290 1768.310 2674.470 ;
        RECT 1767.130 2671.690 1768.310 2672.870 ;
        RECT 1767.130 2493.290 1768.310 2494.470 ;
        RECT 1767.130 2491.690 1768.310 2492.870 ;
        RECT 1767.130 2313.290 1768.310 2314.470 ;
        RECT 1767.130 2311.690 1768.310 2312.870 ;
        RECT 1767.130 2133.290 1768.310 2134.470 ;
        RECT 1767.130 2131.690 1768.310 2132.870 ;
        RECT 1767.130 1953.290 1768.310 1954.470 ;
        RECT 1767.130 1951.690 1768.310 1952.870 ;
        RECT 1767.130 1773.290 1768.310 1774.470 ;
        RECT 1767.130 1771.690 1768.310 1772.870 ;
        RECT 1767.130 1593.290 1768.310 1594.470 ;
        RECT 1767.130 1591.690 1768.310 1592.870 ;
        RECT 1767.130 1413.290 1768.310 1414.470 ;
        RECT 1767.130 1411.690 1768.310 1412.870 ;
        RECT 1767.130 1233.290 1768.310 1234.470 ;
        RECT 1767.130 1231.690 1768.310 1232.870 ;
        RECT 1767.130 1053.290 1768.310 1054.470 ;
        RECT 1767.130 1051.690 1768.310 1052.870 ;
        RECT 1767.130 873.290 1768.310 874.470 ;
        RECT 1767.130 871.690 1768.310 872.870 ;
        RECT 1767.130 693.290 1768.310 694.470 ;
        RECT 1767.130 691.690 1768.310 692.870 ;
        RECT 1767.130 513.290 1768.310 514.470 ;
        RECT 1767.130 511.690 1768.310 512.870 ;
        RECT 1767.130 333.290 1768.310 334.470 ;
        RECT 1767.130 331.690 1768.310 332.870 ;
        RECT 1767.130 153.290 1768.310 154.470 ;
        RECT 1767.130 151.690 1768.310 152.870 ;
        RECT 1767.130 -35.110 1768.310 -33.930 ;
        RECT 1767.130 -36.710 1768.310 -35.530 ;
        RECT 1947.130 3555.210 1948.310 3556.390 ;
        RECT 1947.130 3553.610 1948.310 3554.790 ;
        RECT 1947.130 3393.290 1948.310 3394.470 ;
        RECT 1947.130 3391.690 1948.310 3392.870 ;
        RECT 1947.130 3213.290 1948.310 3214.470 ;
        RECT 1947.130 3211.690 1948.310 3212.870 ;
        RECT 1947.130 3033.290 1948.310 3034.470 ;
        RECT 1947.130 3031.690 1948.310 3032.870 ;
        RECT 1947.130 2853.290 1948.310 2854.470 ;
        RECT 1947.130 2851.690 1948.310 2852.870 ;
        RECT 1947.130 2673.290 1948.310 2674.470 ;
        RECT 1947.130 2671.690 1948.310 2672.870 ;
        RECT 1947.130 2493.290 1948.310 2494.470 ;
        RECT 1947.130 2491.690 1948.310 2492.870 ;
        RECT 1947.130 2313.290 1948.310 2314.470 ;
        RECT 1947.130 2311.690 1948.310 2312.870 ;
        RECT 1947.130 2133.290 1948.310 2134.470 ;
        RECT 1947.130 2131.690 1948.310 2132.870 ;
        RECT 1947.130 1953.290 1948.310 1954.470 ;
        RECT 1947.130 1951.690 1948.310 1952.870 ;
        RECT 1947.130 1773.290 1948.310 1774.470 ;
        RECT 1947.130 1771.690 1948.310 1772.870 ;
        RECT 1947.130 1593.290 1948.310 1594.470 ;
        RECT 1947.130 1591.690 1948.310 1592.870 ;
        RECT 1947.130 1413.290 1948.310 1414.470 ;
        RECT 1947.130 1411.690 1948.310 1412.870 ;
        RECT 1947.130 1233.290 1948.310 1234.470 ;
        RECT 1947.130 1231.690 1948.310 1232.870 ;
        RECT 1947.130 1053.290 1948.310 1054.470 ;
        RECT 1947.130 1051.690 1948.310 1052.870 ;
        RECT 1947.130 873.290 1948.310 874.470 ;
        RECT 1947.130 871.690 1948.310 872.870 ;
        RECT 1947.130 693.290 1948.310 694.470 ;
        RECT 1947.130 691.690 1948.310 692.870 ;
        RECT 1947.130 513.290 1948.310 514.470 ;
        RECT 1947.130 511.690 1948.310 512.870 ;
        RECT 1947.130 333.290 1948.310 334.470 ;
        RECT 1947.130 331.690 1948.310 332.870 ;
        RECT 1947.130 153.290 1948.310 154.470 ;
        RECT 1947.130 151.690 1948.310 152.870 ;
        RECT 1947.130 -35.110 1948.310 -33.930 ;
        RECT 1947.130 -36.710 1948.310 -35.530 ;
        RECT 2127.130 3555.210 2128.310 3556.390 ;
        RECT 2127.130 3553.610 2128.310 3554.790 ;
        RECT 2127.130 3393.290 2128.310 3394.470 ;
        RECT 2127.130 3391.690 2128.310 3392.870 ;
        RECT 2127.130 3213.290 2128.310 3214.470 ;
        RECT 2127.130 3211.690 2128.310 3212.870 ;
        RECT 2127.130 3033.290 2128.310 3034.470 ;
        RECT 2127.130 3031.690 2128.310 3032.870 ;
        RECT 2127.130 2853.290 2128.310 2854.470 ;
        RECT 2127.130 2851.690 2128.310 2852.870 ;
        RECT 2127.130 2673.290 2128.310 2674.470 ;
        RECT 2127.130 2671.690 2128.310 2672.870 ;
        RECT 2127.130 2493.290 2128.310 2494.470 ;
        RECT 2127.130 2491.690 2128.310 2492.870 ;
        RECT 2127.130 2313.290 2128.310 2314.470 ;
        RECT 2127.130 2311.690 2128.310 2312.870 ;
        RECT 2127.130 2133.290 2128.310 2134.470 ;
        RECT 2127.130 2131.690 2128.310 2132.870 ;
        RECT 2127.130 1953.290 2128.310 1954.470 ;
        RECT 2127.130 1951.690 2128.310 1952.870 ;
        RECT 2127.130 1773.290 2128.310 1774.470 ;
        RECT 2127.130 1771.690 2128.310 1772.870 ;
        RECT 2127.130 1593.290 2128.310 1594.470 ;
        RECT 2127.130 1591.690 2128.310 1592.870 ;
        RECT 2127.130 1413.290 2128.310 1414.470 ;
        RECT 2127.130 1411.690 2128.310 1412.870 ;
        RECT 2127.130 1233.290 2128.310 1234.470 ;
        RECT 2127.130 1231.690 2128.310 1232.870 ;
        RECT 2127.130 1053.290 2128.310 1054.470 ;
        RECT 2127.130 1051.690 2128.310 1052.870 ;
        RECT 2127.130 873.290 2128.310 874.470 ;
        RECT 2127.130 871.690 2128.310 872.870 ;
        RECT 2127.130 693.290 2128.310 694.470 ;
        RECT 2127.130 691.690 2128.310 692.870 ;
        RECT 2127.130 513.290 2128.310 514.470 ;
        RECT 2127.130 511.690 2128.310 512.870 ;
        RECT 2127.130 333.290 2128.310 334.470 ;
        RECT 2127.130 331.690 2128.310 332.870 ;
        RECT 2127.130 153.290 2128.310 154.470 ;
        RECT 2127.130 151.690 2128.310 152.870 ;
        RECT 2127.130 -35.110 2128.310 -33.930 ;
        RECT 2127.130 -36.710 2128.310 -35.530 ;
        RECT 2307.130 3555.210 2308.310 3556.390 ;
        RECT 2307.130 3553.610 2308.310 3554.790 ;
        RECT 2307.130 3393.290 2308.310 3394.470 ;
        RECT 2307.130 3391.690 2308.310 3392.870 ;
        RECT 2307.130 3213.290 2308.310 3214.470 ;
        RECT 2307.130 3211.690 2308.310 3212.870 ;
        RECT 2307.130 3033.290 2308.310 3034.470 ;
        RECT 2307.130 3031.690 2308.310 3032.870 ;
        RECT 2307.130 2853.290 2308.310 2854.470 ;
        RECT 2307.130 2851.690 2308.310 2852.870 ;
        RECT 2307.130 2673.290 2308.310 2674.470 ;
        RECT 2307.130 2671.690 2308.310 2672.870 ;
        RECT 2307.130 2493.290 2308.310 2494.470 ;
        RECT 2307.130 2491.690 2308.310 2492.870 ;
        RECT 2307.130 2313.290 2308.310 2314.470 ;
        RECT 2307.130 2311.690 2308.310 2312.870 ;
        RECT 2307.130 2133.290 2308.310 2134.470 ;
        RECT 2307.130 2131.690 2308.310 2132.870 ;
        RECT 2307.130 1953.290 2308.310 1954.470 ;
        RECT 2307.130 1951.690 2308.310 1952.870 ;
        RECT 2307.130 1773.290 2308.310 1774.470 ;
        RECT 2307.130 1771.690 2308.310 1772.870 ;
        RECT 2307.130 1593.290 2308.310 1594.470 ;
        RECT 2307.130 1591.690 2308.310 1592.870 ;
        RECT 2307.130 1413.290 2308.310 1414.470 ;
        RECT 2307.130 1411.690 2308.310 1412.870 ;
        RECT 2307.130 1233.290 2308.310 1234.470 ;
        RECT 2307.130 1231.690 2308.310 1232.870 ;
        RECT 2307.130 1053.290 2308.310 1054.470 ;
        RECT 2307.130 1051.690 2308.310 1052.870 ;
        RECT 2307.130 873.290 2308.310 874.470 ;
        RECT 2307.130 871.690 2308.310 872.870 ;
        RECT 2307.130 693.290 2308.310 694.470 ;
        RECT 2307.130 691.690 2308.310 692.870 ;
        RECT 2307.130 513.290 2308.310 514.470 ;
        RECT 2307.130 511.690 2308.310 512.870 ;
        RECT 2307.130 333.290 2308.310 334.470 ;
        RECT 2307.130 331.690 2308.310 332.870 ;
        RECT 2307.130 153.290 2308.310 154.470 ;
        RECT 2307.130 151.690 2308.310 152.870 ;
        RECT 2307.130 -35.110 2308.310 -33.930 ;
        RECT 2307.130 -36.710 2308.310 -35.530 ;
        RECT 2487.130 3555.210 2488.310 3556.390 ;
        RECT 2487.130 3553.610 2488.310 3554.790 ;
        RECT 2487.130 3393.290 2488.310 3394.470 ;
        RECT 2487.130 3391.690 2488.310 3392.870 ;
        RECT 2487.130 3213.290 2488.310 3214.470 ;
        RECT 2487.130 3211.690 2488.310 3212.870 ;
        RECT 2487.130 3033.290 2488.310 3034.470 ;
        RECT 2487.130 3031.690 2488.310 3032.870 ;
        RECT 2487.130 2853.290 2488.310 2854.470 ;
        RECT 2487.130 2851.690 2488.310 2852.870 ;
        RECT 2487.130 2673.290 2488.310 2674.470 ;
        RECT 2487.130 2671.690 2488.310 2672.870 ;
        RECT 2487.130 2493.290 2488.310 2494.470 ;
        RECT 2487.130 2491.690 2488.310 2492.870 ;
        RECT 2487.130 2313.290 2488.310 2314.470 ;
        RECT 2487.130 2311.690 2488.310 2312.870 ;
        RECT 2487.130 2133.290 2488.310 2134.470 ;
        RECT 2487.130 2131.690 2488.310 2132.870 ;
        RECT 2487.130 1953.290 2488.310 1954.470 ;
        RECT 2487.130 1951.690 2488.310 1952.870 ;
        RECT 2487.130 1773.290 2488.310 1774.470 ;
        RECT 2487.130 1771.690 2488.310 1772.870 ;
        RECT 2487.130 1593.290 2488.310 1594.470 ;
        RECT 2487.130 1591.690 2488.310 1592.870 ;
        RECT 2487.130 1413.290 2488.310 1414.470 ;
        RECT 2487.130 1411.690 2488.310 1412.870 ;
        RECT 2487.130 1233.290 2488.310 1234.470 ;
        RECT 2487.130 1231.690 2488.310 1232.870 ;
        RECT 2487.130 1053.290 2488.310 1054.470 ;
        RECT 2487.130 1051.690 2488.310 1052.870 ;
        RECT 2487.130 873.290 2488.310 874.470 ;
        RECT 2487.130 871.690 2488.310 872.870 ;
        RECT 2487.130 693.290 2488.310 694.470 ;
        RECT 2487.130 691.690 2488.310 692.870 ;
        RECT 2487.130 513.290 2488.310 514.470 ;
        RECT 2487.130 511.690 2488.310 512.870 ;
        RECT 2487.130 333.290 2488.310 334.470 ;
        RECT 2487.130 331.690 2488.310 332.870 ;
        RECT 2487.130 153.290 2488.310 154.470 ;
        RECT 2487.130 151.690 2488.310 152.870 ;
        RECT 2487.130 -35.110 2488.310 -33.930 ;
        RECT 2487.130 -36.710 2488.310 -35.530 ;
        RECT 2667.130 3555.210 2668.310 3556.390 ;
        RECT 2667.130 3553.610 2668.310 3554.790 ;
        RECT 2667.130 3393.290 2668.310 3394.470 ;
        RECT 2667.130 3391.690 2668.310 3392.870 ;
        RECT 2667.130 3213.290 2668.310 3214.470 ;
        RECT 2667.130 3211.690 2668.310 3212.870 ;
        RECT 2667.130 3033.290 2668.310 3034.470 ;
        RECT 2667.130 3031.690 2668.310 3032.870 ;
        RECT 2667.130 2853.290 2668.310 2854.470 ;
        RECT 2667.130 2851.690 2668.310 2852.870 ;
        RECT 2667.130 2673.290 2668.310 2674.470 ;
        RECT 2667.130 2671.690 2668.310 2672.870 ;
        RECT 2667.130 2493.290 2668.310 2494.470 ;
        RECT 2667.130 2491.690 2668.310 2492.870 ;
        RECT 2667.130 2313.290 2668.310 2314.470 ;
        RECT 2667.130 2311.690 2668.310 2312.870 ;
        RECT 2667.130 2133.290 2668.310 2134.470 ;
        RECT 2667.130 2131.690 2668.310 2132.870 ;
        RECT 2667.130 1953.290 2668.310 1954.470 ;
        RECT 2667.130 1951.690 2668.310 1952.870 ;
        RECT 2667.130 1773.290 2668.310 1774.470 ;
        RECT 2667.130 1771.690 2668.310 1772.870 ;
        RECT 2667.130 1593.290 2668.310 1594.470 ;
        RECT 2667.130 1591.690 2668.310 1592.870 ;
        RECT 2667.130 1413.290 2668.310 1414.470 ;
        RECT 2667.130 1411.690 2668.310 1412.870 ;
        RECT 2667.130 1233.290 2668.310 1234.470 ;
        RECT 2667.130 1231.690 2668.310 1232.870 ;
        RECT 2667.130 1053.290 2668.310 1054.470 ;
        RECT 2667.130 1051.690 2668.310 1052.870 ;
        RECT 2667.130 873.290 2668.310 874.470 ;
        RECT 2667.130 871.690 2668.310 872.870 ;
        RECT 2667.130 693.290 2668.310 694.470 ;
        RECT 2667.130 691.690 2668.310 692.870 ;
        RECT 2667.130 513.290 2668.310 514.470 ;
        RECT 2667.130 511.690 2668.310 512.870 ;
        RECT 2667.130 333.290 2668.310 334.470 ;
        RECT 2667.130 331.690 2668.310 332.870 ;
        RECT 2667.130 153.290 2668.310 154.470 ;
        RECT 2667.130 151.690 2668.310 152.870 ;
        RECT 2667.130 -35.110 2668.310 -33.930 ;
        RECT 2667.130 -36.710 2668.310 -35.530 ;
        RECT 2847.130 3555.210 2848.310 3556.390 ;
        RECT 2847.130 3553.610 2848.310 3554.790 ;
        RECT 2847.130 3393.290 2848.310 3394.470 ;
        RECT 2847.130 3391.690 2848.310 3392.870 ;
        RECT 2847.130 3213.290 2848.310 3214.470 ;
        RECT 2847.130 3211.690 2848.310 3212.870 ;
        RECT 2847.130 3033.290 2848.310 3034.470 ;
        RECT 2847.130 3031.690 2848.310 3032.870 ;
        RECT 2847.130 2853.290 2848.310 2854.470 ;
        RECT 2847.130 2851.690 2848.310 2852.870 ;
        RECT 2847.130 2673.290 2848.310 2674.470 ;
        RECT 2847.130 2671.690 2848.310 2672.870 ;
        RECT 2847.130 2493.290 2848.310 2494.470 ;
        RECT 2847.130 2491.690 2848.310 2492.870 ;
        RECT 2847.130 2313.290 2848.310 2314.470 ;
        RECT 2847.130 2311.690 2848.310 2312.870 ;
        RECT 2847.130 2133.290 2848.310 2134.470 ;
        RECT 2847.130 2131.690 2848.310 2132.870 ;
        RECT 2847.130 1953.290 2848.310 1954.470 ;
        RECT 2847.130 1951.690 2848.310 1952.870 ;
        RECT 2847.130 1773.290 2848.310 1774.470 ;
        RECT 2847.130 1771.690 2848.310 1772.870 ;
        RECT 2847.130 1593.290 2848.310 1594.470 ;
        RECT 2847.130 1591.690 2848.310 1592.870 ;
        RECT 2847.130 1413.290 2848.310 1414.470 ;
        RECT 2847.130 1411.690 2848.310 1412.870 ;
        RECT 2847.130 1233.290 2848.310 1234.470 ;
        RECT 2847.130 1231.690 2848.310 1232.870 ;
        RECT 2847.130 1053.290 2848.310 1054.470 ;
        RECT 2847.130 1051.690 2848.310 1052.870 ;
        RECT 2847.130 873.290 2848.310 874.470 ;
        RECT 2847.130 871.690 2848.310 872.870 ;
        RECT 2847.130 693.290 2848.310 694.470 ;
        RECT 2847.130 691.690 2848.310 692.870 ;
        RECT 2847.130 513.290 2848.310 514.470 ;
        RECT 2847.130 511.690 2848.310 512.870 ;
        RECT 2847.130 333.290 2848.310 334.470 ;
        RECT 2847.130 331.690 2848.310 332.870 ;
        RECT 2847.130 153.290 2848.310 154.470 ;
        RECT 2847.130 151.690 2848.310 152.870 ;
        RECT 2847.130 -35.110 2848.310 -33.930 ;
        RECT 2847.130 -36.710 2848.310 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3393.290 2960.890 3394.470 ;
        RECT 2959.710 3391.690 2960.890 3392.870 ;
        RECT 2959.710 3213.290 2960.890 3214.470 ;
        RECT 2959.710 3211.690 2960.890 3212.870 ;
        RECT 2959.710 3033.290 2960.890 3034.470 ;
        RECT 2959.710 3031.690 2960.890 3032.870 ;
        RECT 2959.710 2853.290 2960.890 2854.470 ;
        RECT 2959.710 2851.690 2960.890 2852.870 ;
        RECT 2959.710 2673.290 2960.890 2674.470 ;
        RECT 2959.710 2671.690 2960.890 2672.870 ;
        RECT 2959.710 2493.290 2960.890 2494.470 ;
        RECT 2959.710 2491.690 2960.890 2492.870 ;
        RECT 2959.710 2313.290 2960.890 2314.470 ;
        RECT 2959.710 2311.690 2960.890 2312.870 ;
        RECT 2959.710 2133.290 2960.890 2134.470 ;
        RECT 2959.710 2131.690 2960.890 2132.870 ;
        RECT 2959.710 1953.290 2960.890 1954.470 ;
        RECT 2959.710 1951.690 2960.890 1952.870 ;
        RECT 2959.710 1773.290 2960.890 1774.470 ;
        RECT 2959.710 1771.690 2960.890 1772.870 ;
        RECT 2959.710 1593.290 2960.890 1594.470 ;
        RECT 2959.710 1591.690 2960.890 1592.870 ;
        RECT 2959.710 1413.290 2960.890 1414.470 ;
        RECT 2959.710 1411.690 2960.890 1412.870 ;
        RECT 2959.710 1233.290 2960.890 1234.470 ;
        RECT 2959.710 1231.690 2960.890 1232.870 ;
        RECT 2959.710 1053.290 2960.890 1054.470 ;
        RECT 2959.710 1051.690 2960.890 1052.870 ;
        RECT 2959.710 873.290 2960.890 874.470 ;
        RECT 2959.710 871.690 2960.890 872.870 ;
        RECT 2959.710 693.290 2960.890 694.470 ;
        RECT 2959.710 691.690 2960.890 692.870 ;
        RECT 2959.710 513.290 2960.890 514.470 ;
        RECT 2959.710 511.690 2960.890 512.870 ;
        RECT 2959.710 333.290 2960.890 334.470 ;
        RECT 2959.710 331.690 2960.890 332.870 ;
        RECT 2959.710 153.290 2960.890 154.470 ;
        RECT 2959.710 151.690 2960.890 152.870 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.130 3556.450 -39.230 3556.510 ;
        RECT 146.270 3556.450 149.170 3556.510 ;
        RECT 326.270 3556.450 329.170 3556.510 ;
        RECT 506.270 3556.450 509.170 3556.510 ;
        RECT 686.270 3556.450 689.170 3556.510 ;
        RECT 866.270 3556.450 869.170 3556.510 ;
        RECT 1046.270 3556.450 1049.170 3556.510 ;
        RECT 1226.270 3556.450 1229.170 3556.510 ;
        RECT 1406.270 3556.450 1409.170 3556.510 ;
        RECT 1586.270 3556.450 1589.170 3556.510 ;
        RECT 1766.270 3556.450 1769.170 3556.510 ;
        RECT 1946.270 3556.450 1949.170 3556.510 ;
        RECT 2126.270 3556.450 2129.170 3556.510 ;
        RECT 2306.270 3556.450 2309.170 3556.510 ;
        RECT 2486.270 3556.450 2489.170 3556.510 ;
        RECT 2666.270 3556.450 2669.170 3556.510 ;
        RECT 2846.270 3556.450 2849.170 3556.510 ;
        RECT 2958.850 3556.450 2961.750 3556.510 ;
        RECT -42.130 3553.550 2961.750 3556.450 ;
        RECT -42.130 3553.490 -39.230 3553.550 ;
        RECT 146.270 3553.490 149.170 3553.550 ;
        RECT 326.270 3553.490 329.170 3553.550 ;
        RECT 506.270 3553.490 509.170 3553.550 ;
        RECT 686.270 3553.490 689.170 3553.550 ;
        RECT 866.270 3553.490 869.170 3553.550 ;
        RECT 1046.270 3553.490 1049.170 3553.550 ;
        RECT 1226.270 3553.490 1229.170 3553.550 ;
        RECT 1406.270 3553.490 1409.170 3553.550 ;
        RECT 1586.270 3553.490 1589.170 3553.550 ;
        RECT 1766.270 3553.490 1769.170 3553.550 ;
        RECT 1946.270 3553.490 1949.170 3553.550 ;
        RECT 2126.270 3553.490 2129.170 3553.550 ;
        RECT 2306.270 3553.490 2309.170 3553.550 ;
        RECT 2486.270 3553.490 2489.170 3553.550 ;
        RECT 2666.270 3553.490 2669.170 3553.550 ;
        RECT 2846.270 3553.490 2849.170 3553.550 ;
        RECT 2958.850 3553.490 2961.750 3553.550 ;
        RECT -42.130 3394.530 -39.230 3394.590 ;
        RECT 146.270 3394.530 149.170 3394.590 ;
        RECT 326.270 3394.530 329.170 3394.590 ;
        RECT 506.270 3394.530 509.170 3394.590 ;
        RECT 686.270 3394.530 689.170 3394.590 ;
        RECT 866.270 3394.530 869.170 3394.590 ;
        RECT 1046.270 3394.530 1049.170 3394.590 ;
        RECT 1226.270 3394.530 1229.170 3394.590 ;
        RECT 1406.270 3394.530 1409.170 3394.590 ;
        RECT 1586.270 3394.530 1589.170 3394.590 ;
        RECT 1766.270 3394.530 1769.170 3394.590 ;
        RECT 1946.270 3394.530 1949.170 3394.590 ;
        RECT 2126.270 3394.530 2129.170 3394.590 ;
        RECT 2306.270 3394.530 2309.170 3394.590 ;
        RECT 2486.270 3394.530 2489.170 3394.590 ;
        RECT 2666.270 3394.530 2669.170 3394.590 ;
        RECT 2846.270 3394.530 2849.170 3394.590 ;
        RECT 2958.850 3394.530 2961.750 3394.590 ;
        RECT -42.130 3391.630 2961.750 3394.530 ;
        RECT -42.130 3391.570 -39.230 3391.630 ;
        RECT 146.270 3391.570 149.170 3391.630 ;
        RECT 326.270 3391.570 329.170 3391.630 ;
        RECT 506.270 3391.570 509.170 3391.630 ;
        RECT 686.270 3391.570 689.170 3391.630 ;
        RECT 866.270 3391.570 869.170 3391.630 ;
        RECT 1046.270 3391.570 1049.170 3391.630 ;
        RECT 1226.270 3391.570 1229.170 3391.630 ;
        RECT 1406.270 3391.570 1409.170 3391.630 ;
        RECT 1586.270 3391.570 1589.170 3391.630 ;
        RECT 1766.270 3391.570 1769.170 3391.630 ;
        RECT 1946.270 3391.570 1949.170 3391.630 ;
        RECT 2126.270 3391.570 2129.170 3391.630 ;
        RECT 2306.270 3391.570 2309.170 3391.630 ;
        RECT 2486.270 3391.570 2489.170 3391.630 ;
        RECT 2666.270 3391.570 2669.170 3391.630 ;
        RECT 2846.270 3391.570 2849.170 3391.630 ;
        RECT 2958.850 3391.570 2961.750 3391.630 ;
        RECT -42.130 3214.530 -39.230 3214.590 ;
        RECT 146.270 3214.530 149.170 3214.590 ;
        RECT 326.270 3214.530 329.170 3214.590 ;
        RECT 506.270 3214.530 509.170 3214.590 ;
        RECT 686.270 3214.530 689.170 3214.590 ;
        RECT 866.270 3214.530 869.170 3214.590 ;
        RECT 1046.270 3214.530 1049.170 3214.590 ;
        RECT 1226.270 3214.530 1229.170 3214.590 ;
        RECT 1406.270 3214.530 1409.170 3214.590 ;
        RECT 1586.270 3214.530 1589.170 3214.590 ;
        RECT 1766.270 3214.530 1769.170 3214.590 ;
        RECT 1946.270 3214.530 1949.170 3214.590 ;
        RECT 2126.270 3214.530 2129.170 3214.590 ;
        RECT 2306.270 3214.530 2309.170 3214.590 ;
        RECT 2486.270 3214.530 2489.170 3214.590 ;
        RECT 2666.270 3214.530 2669.170 3214.590 ;
        RECT 2846.270 3214.530 2849.170 3214.590 ;
        RECT 2958.850 3214.530 2961.750 3214.590 ;
        RECT -42.130 3211.630 2961.750 3214.530 ;
        RECT -42.130 3211.570 -39.230 3211.630 ;
        RECT 146.270 3211.570 149.170 3211.630 ;
        RECT 326.270 3211.570 329.170 3211.630 ;
        RECT 506.270 3211.570 509.170 3211.630 ;
        RECT 686.270 3211.570 689.170 3211.630 ;
        RECT 866.270 3211.570 869.170 3211.630 ;
        RECT 1046.270 3211.570 1049.170 3211.630 ;
        RECT 1226.270 3211.570 1229.170 3211.630 ;
        RECT 1406.270 3211.570 1409.170 3211.630 ;
        RECT 1586.270 3211.570 1589.170 3211.630 ;
        RECT 1766.270 3211.570 1769.170 3211.630 ;
        RECT 1946.270 3211.570 1949.170 3211.630 ;
        RECT 2126.270 3211.570 2129.170 3211.630 ;
        RECT 2306.270 3211.570 2309.170 3211.630 ;
        RECT 2486.270 3211.570 2489.170 3211.630 ;
        RECT 2666.270 3211.570 2669.170 3211.630 ;
        RECT 2846.270 3211.570 2849.170 3211.630 ;
        RECT 2958.850 3211.570 2961.750 3211.630 ;
        RECT -42.130 3034.530 -39.230 3034.590 ;
        RECT 146.270 3034.530 149.170 3034.590 ;
        RECT 326.270 3034.530 329.170 3034.590 ;
        RECT 506.270 3034.530 509.170 3034.590 ;
        RECT 686.270 3034.530 689.170 3034.590 ;
        RECT 866.270 3034.530 869.170 3034.590 ;
        RECT 1046.270 3034.530 1049.170 3034.590 ;
        RECT 1226.270 3034.530 1229.170 3034.590 ;
        RECT 1406.270 3034.530 1409.170 3034.590 ;
        RECT 1586.270 3034.530 1589.170 3034.590 ;
        RECT 1766.270 3034.530 1769.170 3034.590 ;
        RECT 1946.270 3034.530 1949.170 3034.590 ;
        RECT 2126.270 3034.530 2129.170 3034.590 ;
        RECT 2306.270 3034.530 2309.170 3034.590 ;
        RECT 2486.270 3034.530 2489.170 3034.590 ;
        RECT 2666.270 3034.530 2669.170 3034.590 ;
        RECT 2846.270 3034.530 2849.170 3034.590 ;
        RECT 2958.850 3034.530 2961.750 3034.590 ;
        RECT -42.130 3031.630 2961.750 3034.530 ;
        RECT -42.130 3031.570 -39.230 3031.630 ;
        RECT 146.270 3031.570 149.170 3031.630 ;
        RECT 326.270 3031.570 329.170 3031.630 ;
        RECT 506.270 3031.570 509.170 3031.630 ;
        RECT 686.270 3031.570 689.170 3031.630 ;
        RECT 866.270 3031.570 869.170 3031.630 ;
        RECT 1046.270 3031.570 1049.170 3031.630 ;
        RECT 1226.270 3031.570 1229.170 3031.630 ;
        RECT 1406.270 3031.570 1409.170 3031.630 ;
        RECT 1586.270 3031.570 1589.170 3031.630 ;
        RECT 1766.270 3031.570 1769.170 3031.630 ;
        RECT 1946.270 3031.570 1949.170 3031.630 ;
        RECT 2126.270 3031.570 2129.170 3031.630 ;
        RECT 2306.270 3031.570 2309.170 3031.630 ;
        RECT 2486.270 3031.570 2489.170 3031.630 ;
        RECT 2666.270 3031.570 2669.170 3031.630 ;
        RECT 2846.270 3031.570 2849.170 3031.630 ;
        RECT 2958.850 3031.570 2961.750 3031.630 ;
        RECT -42.130 2854.530 -39.230 2854.590 ;
        RECT 146.270 2854.530 149.170 2854.590 ;
        RECT 326.270 2854.530 329.170 2854.590 ;
        RECT 506.270 2854.530 509.170 2854.590 ;
        RECT 686.270 2854.530 689.170 2854.590 ;
        RECT 866.270 2854.530 869.170 2854.590 ;
        RECT 1046.270 2854.530 1049.170 2854.590 ;
        RECT 1226.270 2854.530 1229.170 2854.590 ;
        RECT 1406.270 2854.530 1409.170 2854.590 ;
        RECT 1586.270 2854.530 1589.170 2854.590 ;
        RECT 1766.270 2854.530 1769.170 2854.590 ;
        RECT 1946.270 2854.530 1949.170 2854.590 ;
        RECT 2126.270 2854.530 2129.170 2854.590 ;
        RECT 2306.270 2854.530 2309.170 2854.590 ;
        RECT 2486.270 2854.530 2489.170 2854.590 ;
        RECT 2666.270 2854.530 2669.170 2854.590 ;
        RECT 2846.270 2854.530 2849.170 2854.590 ;
        RECT 2958.850 2854.530 2961.750 2854.590 ;
        RECT -42.130 2851.630 2961.750 2854.530 ;
        RECT -42.130 2851.570 -39.230 2851.630 ;
        RECT 146.270 2851.570 149.170 2851.630 ;
        RECT 326.270 2851.570 329.170 2851.630 ;
        RECT 506.270 2851.570 509.170 2851.630 ;
        RECT 686.270 2851.570 689.170 2851.630 ;
        RECT 866.270 2851.570 869.170 2851.630 ;
        RECT 1046.270 2851.570 1049.170 2851.630 ;
        RECT 1226.270 2851.570 1229.170 2851.630 ;
        RECT 1406.270 2851.570 1409.170 2851.630 ;
        RECT 1586.270 2851.570 1589.170 2851.630 ;
        RECT 1766.270 2851.570 1769.170 2851.630 ;
        RECT 1946.270 2851.570 1949.170 2851.630 ;
        RECT 2126.270 2851.570 2129.170 2851.630 ;
        RECT 2306.270 2851.570 2309.170 2851.630 ;
        RECT 2486.270 2851.570 2489.170 2851.630 ;
        RECT 2666.270 2851.570 2669.170 2851.630 ;
        RECT 2846.270 2851.570 2849.170 2851.630 ;
        RECT 2958.850 2851.570 2961.750 2851.630 ;
        RECT -42.130 2674.530 -39.230 2674.590 ;
        RECT 146.270 2674.530 149.170 2674.590 ;
        RECT 326.270 2674.530 329.170 2674.590 ;
        RECT 506.270 2674.530 509.170 2674.590 ;
        RECT 686.270 2674.530 689.170 2674.590 ;
        RECT 866.270 2674.530 869.170 2674.590 ;
        RECT 1046.270 2674.530 1049.170 2674.590 ;
        RECT 1226.270 2674.530 1229.170 2674.590 ;
        RECT 1406.270 2674.530 1409.170 2674.590 ;
        RECT 1586.270 2674.530 1589.170 2674.590 ;
        RECT 1766.270 2674.530 1769.170 2674.590 ;
        RECT 1946.270 2674.530 1949.170 2674.590 ;
        RECT 2126.270 2674.530 2129.170 2674.590 ;
        RECT 2306.270 2674.530 2309.170 2674.590 ;
        RECT 2486.270 2674.530 2489.170 2674.590 ;
        RECT 2666.270 2674.530 2669.170 2674.590 ;
        RECT 2846.270 2674.530 2849.170 2674.590 ;
        RECT 2958.850 2674.530 2961.750 2674.590 ;
        RECT -42.130 2671.630 2961.750 2674.530 ;
        RECT -42.130 2671.570 -39.230 2671.630 ;
        RECT 146.270 2671.570 149.170 2671.630 ;
        RECT 326.270 2671.570 329.170 2671.630 ;
        RECT 506.270 2671.570 509.170 2671.630 ;
        RECT 686.270 2671.570 689.170 2671.630 ;
        RECT 866.270 2671.570 869.170 2671.630 ;
        RECT 1046.270 2671.570 1049.170 2671.630 ;
        RECT 1226.270 2671.570 1229.170 2671.630 ;
        RECT 1406.270 2671.570 1409.170 2671.630 ;
        RECT 1586.270 2671.570 1589.170 2671.630 ;
        RECT 1766.270 2671.570 1769.170 2671.630 ;
        RECT 1946.270 2671.570 1949.170 2671.630 ;
        RECT 2126.270 2671.570 2129.170 2671.630 ;
        RECT 2306.270 2671.570 2309.170 2671.630 ;
        RECT 2486.270 2671.570 2489.170 2671.630 ;
        RECT 2666.270 2671.570 2669.170 2671.630 ;
        RECT 2846.270 2671.570 2849.170 2671.630 ;
        RECT 2958.850 2671.570 2961.750 2671.630 ;
        RECT -42.130 2494.530 -39.230 2494.590 ;
        RECT 146.270 2494.530 149.170 2494.590 ;
        RECT 326.270 2494.530 329.170 2494.590 ;
        RECT 506.270 2494.530 509.170 2494.590 ;
        RECT 686.270 2494.530 689.170 2494.590 ;
        RECT 866.270 2494.530 869.170 2494.590 ;
        RECT 1046.270 2494.530 1049.170 2494.590 ;
        RECT 1226.270 2494.530 1229.170 2494.590 ;
        RECT 1406.270 2494.530 1409.170 2494.590 ;
        RECT 1586.270 2494.530 1589.170 2494.590 ;
        RECT 1766.270 2494.530 1769.170 2494.590 ;
        RECT 1946.270 2494.530 1949.170 2494.590 ;
        RECT 2126.270 2494.530 2129.170 2494.590 ;
        RECT 2306.270 2494.530 2309.170 2494.590 ;
        RECT 2486.270 2494.530 2489.170 2494.590 ;
        RECT 2666.270 2494.530 2669.170 2494.590 ;
        RECT 2846.270 2494.530 2849.170 2494.590 ;
        RECT 2958.850 2494.530 2961.750 2494.590 ;
        RECT -42.130 2491.630 2961.750 2494.530 ;
        RECT -42.130 2491.570 -39.230 2491.630 ;
        RECT 146.270 2491.570 149.170 2491.630 ;
        RECT 326.270 2491.570 329.170 2491.630 ;
        RECT 506.270 2491.570 509.170 2491.630 ;
        RECT 686.270 2491.570 689.170 2491.630 ;
        RECT 866.270 2491.570 869.170 2491.630 ;
        RECT 1046.270 2491.570 1049.170 2491.630 ;
        RECT 1226.270 2491.570 1229.170 2491.630 ;
        RECT 1406.270 2491.570 1409.170 2491.630 ;
        RECT 1586.270 2491.570 1589.170 2491.630 ;
        RECT 1766.270 2491.570 1769.170 2491.630 ;
        RECT 1946.270 2491.570 1949.170 2491.630 ;
        RECT 2126.270 2491.570 2129.170 2491.630 ;
        RECT 2306.270 2491.570 2309.170 2491.630 ;
        RECT 2486.270 2491.570 2489.170 2491.630 ;
        RECT 2666.270 2491.570 2669.170 2491.630 ;
        RECT 2846.270 2491.570 2849.170 2491.630 ;
        RECT 2958.850 2491.570 2961.750 2491.630 ;
        RECT -42.130 2314.530 -39.230 2314.590 ;
        RECT 146.270 2314.530 149.170 2314.590 ;
        RECT 326.270 2314.530 329.170 2314.590 ;
        RECT 506.270 2314.530 509.170 2314.590 ;
        RECT 686.270 2314.530 689.170 2314.590 ;
        RECT 866.270 2314.530 869.170 2314.590 ;
        RECT 1046.270 2314.530 1049.170 2314.590 ;
        RECT 1226.270 2314.530 1229.170 2314.590 ;
        RECT 1406.270 2314.530 1409.170 2314.590 ;
        RECT 1586.270 2314.530 1589.170 2314.590 ;
        RECT 1766.270 2314.530 1769.170 2314.590 ;
        RECT 1946.270 2314.530 1949.170 2314.590 ;
        RECT 2126.270 2314.530 2129.170 2314.590 ;
        RECT 2306.270 2314.530 2309.170 2314.590 ;
        RECT 2486.270 2314.530 2489.170 2314.590 ;
        RECT 2666.270 2314.530 2669.170 2314.590 ;
        RECT 2846.270 2314.530 2849.170 2314.590 ;
        RECT 2958.850 2314.530 2961.750 2314.590 ;
        RECT -42.130 2311.630 2961.750 2314.530 ;
        RECT -42.130 2311.570 -39.230 2311.630 ;
        RECT 146.270 2311.570 149.170 2311.630 ;
        RECT 326.270 2311.570 329.170 2311.630 ;
        RECT 506.270 2311.570 509.170 2311.630 ;
        RECT 686.270 2311.570 689.170 2311.630 ;
        RECT 866.270 2311.570 869.170 2311.630 ;
        RECT 1046.270 2311.570 1049.170 2311.630 ;
        RECT 1226.270 2311.570 1229.170 2311.630 ;
        RECT 1406.270 2311.570 1409.170 2311.630 ;
        RECT 1586.270 2311.570 1589.170 2311.630 ;
        RECT 1766.270 2311.570 1769.170 2311.630 ;
        RECT 1946.270 2311.570 1949.170 2311.630 ;
        RECT 2126.270 2311.570 2129.170 2311.630 ;
        RECT 2306.270 2311.570 2309.170 2311.630 ;
        RECT 2486.270 2311.570 2489.170 2311.630 ;
        RECT 2666.270 2311.570 2669.170 2311.630 ;
        RECT 2846.270 2311.570 2849.170 2311.630 ;
        RECT 2958.850 2311.570 2961.750 2311.630 ;
        RECT -42.130 2134.530 -39.230 2134.590 ;
        RECT 146.270 2134.530 149.170 2134.590 ;
        RECT 326.270 2134.530 329.170 2134.590 ;
        RECT 506.270 2134.530 509.170 2134.590 ;
        RECT 686.270 2134.530 689.170 2134.590 ;
        RECT 866.270 2134.530 869.170 2134.590 ;
        RECT 1046.270 2134.530 1049.170 2134.590 ;
        RECT 1226.270 2134.530 1229.170 2134.590 ;
        RECT 1406.270 2134.530 1409.170 2134.590 ;
        RECT 1586.270 2134.530 1589.170 2134.590 ;
        RECT 1766.270 2134.530 1769.170 2134.590 ;
        RECT 1946.270 2134.530 1949.170 2134.590 ;
        RECT 2126.270 2134.530 2129.170 2134.590 ;
        RECT 2306.270 2134.530 2309.170 2134.590 ;
        RECT 2486.270 2134.530 2489.170 2134.590 ;
        RECT 2666.270 2134.530 2669.170 2134.590 ;
        RECT 2846.270 2134.530 2849.170 2134.590 ;
        RECT 2958.850 2134.530 2961.750 2134.590 ;
        RECT -42.130 2131.630 2961.750 2134.530 ;
        RECT -42.130 2131.570 -39.230 2131.630 ;
        RECT 146.270 2131.570 149.170 2131.630 ;
        RECT 326.270 2131.570 329.170 2131.630 ;
        RECT 506.270 2131.570 509.170 2131.630 ;
        RECT 686.270 2131.570 689.170 2131.630 ;
        RECT 866.270 2131.570 869.170 2131.630 ;
        RECT 1046.270 2131.570 1049.170 2131.630 ;
        RECT 1226.270 2131.570 1229.170 2131.630 ;
        RECT 1406.270 2131.570 1409.170 2131.630 ;
        RECT 1586.270 2131.570 1589.170 2131.630 ;
        RECT 1766.270 2131.570 1769.170 2131.630 ;
        RECT 1946.270 2131.570 1949.170 2131.630 ;
        RECT 2126.270 2131.570 2129.170 2131.630 ;
        RECT 2306.270 2131.570 2309.170 2131.630 ;
        RECT 2486.270 2131.570 2489.170 2131.630 ;
        RECT 2666.270 2131.570 2669.170 2131.630 ;
        RECT 2846.270 2131.570 2849.170 2131.630 ;
        RECT 2958.850 2131.570 2961.750 2131.630 ;
        RECT -42.130 1954.530 -39.230 1954.590 ;
        RECT 146.270 1954.530 149.170 1954.590 ;
        RECT 326.270 1954.530 329.170 1954.590 ;
        RECT 506.270 1954.530 509.170 1954.590 ;
        RECT 686.270 1954.530 689.170 1954.590 ;
        RECT 866.270 1954.530 869.170 1954.590 ;
        RECT 1046.270 1954.530 1049.170 1954.590 ;
        RECT 1226.270 1954.530 1229.170 1954.590 ;
        RECT 1406.270 1954.530 1409.170 1954.590 ;
        RECT 1586.270 1954.530 1589.170 1954.590 ;
        RECT 1766.270 1954.530 1769.170 1954.590 ;
        RECT 1946.270 1954.530 1949.170 1954.590 ;
        RECT 2126.270 1954.530 2129.170 1954.590 ;
        RECT 2306.270 1954.530 2309.170 1954.590 ;
        RECT 2486.270 1954.530 2489.170 1954.590 ;
        RECT 2666.270 1954.530 2669.170 1954.590 ;
        RECT 2846.270 1954.530 2849.170 1954.590 ;
        RECT 2958.850 1954.530 2961.750 1954.590 ;
        RECT -42.130 1951.630 2961.750 1954.530 ;
        RECT -42.130 1951.570 -39.230 1951.630 ;
        RECT 146.270 1951.570 149.170 1951.630 ;
        RECT 326.270 1951.570 329.170 1951.630 ;
        RECT 506.270 1951.570 509.170 1951.630 ;
        RECT 686.270 1951.570 689.170 1951.630 ;
        RECT 866.270 1951.570 869.170 1951.630 ;
        RECT 1046.270 1951.570 1049.170 1951.630 ;
        RECT 1226.270 1951.570 1229.170 1951.630 ;
        RECT 1406.270 1951.570 1409.170 1951.630 ;
        RECT 1586.270 1951.570 1589.170 1951.630 ;
        RECT 1766.270 1951.570 1769.170 1951.630 ;
        RECT 1946.270 1951.570 1949.170 1951.630 ;
        RECT 2126.270 1951.570 2129.170 1951.630 ;
        RECT 2306.270 1951.570 2309.170 1951.630 ;
        RECT 2486.270 1951.570 2489.170 1951.630 ;
        RECT 2666.270 1951.570 2669.170 1951.630 ;
        RECT 2846.270 1951.570 2849.170 1951.630 ;
        RECT 2958.850 1951.570 2961.750 1951.630 ;
        RECT -42.130 1774.530 -39.230 1774.590 ;
        RECT 146.270 1774.530 149.170 1774.590 ;
        RECT 326.270 1774.530 329.170 1774.590 ;
        RECT 506.270 1774.530 509.170 1774.590 ;
        RECT 686.270 1774.530 689.170 1774.590 ;
        RECT 866.270 1774.530 869.170 1774.590 ;
        RECT 1046.270 1774.530 1049.170 1774.590 ;
        RECT 1226.270 1774.530 1229.170 1774.590 ;
        RECT 1406.270 1774.530 1409.170 1774.590 ;
        RECT 1586.270 1774.530 1589.170 1774.590 ;
        RECT 1766.270 1774.530 1769.170 1774.590 ;
        RECT 1946.270 1774.530 1949.170 1774.590 ;
        RECT 2126.270 1774.530 2129.170 1774.590 ;
        RECT 2306.270 1774.530 2309.170 1774.590 ;
        RECT 2486.270 1774.530 2489.170 1774.590 ;
        RECT 2666.270 1774.530 2669.170 1774.590 ;
        RECT 2846.270 1774.530 2849.170 1774.590 ;
        RECT 2958.850 1774.530 2961.750 1774.590 ;
        RECT -42.130 1771.630 2961.750 1774.530 ;
        RECT -42.130 1771.570 -39.230 1771.630 ;
        RECT 146.270 1771.570 149.170 1771.630 ;
        RECT 326.270 1771.570 329.170 1771.630 ;
        RECT 506.270 1771.570 509.170 1771.630 ;
        RECT 686.270 1771.570 689.170 1771.630 ;
        RECT 866.270 1771.570 869.170 1771.630 ;
        RECT 1046.270 1771.570 1049.170 1771.630 ;
        RECT 1226.270 1771.570 1229.170 1771.630 ;
        RECT 1406.270 1771.570 1409.170 1771.630 ;
        RECT 1586.270 1771.570 1589.170 1771.630 ;
        RECT 1766.270 1771.570 1769.170 1771.630 ;
        RECT 1946.270 1771.570 1949.170 1771.630 ;
        RECT 2126.270 1771.570 2129.170 1771.630 ;
        RECT 2306.270 1771.570 2309.170 1771.630 ;
        RECT 2486.270 1771.570 2489.170 1771.630 ;
        RECT 2666.270 1771.570 2669.170 1771.630 ;
        RECT 2846.270 1771.570 2849.170 1771.630 ;
        RECT 2958.850 1771.570 2961.750 1771.630 ;
        RECT -42.130 1594.530 -39.230 1594.590 ;
        RECT 146.270 1594.530 149.170 1594.590 ;
        RECT 326.270 1594.530 329.170 1594.590 ;
        RECT 506.270 1594.530 509.170 1594.590 ;
        RECT 686.270 1594.530 689.170 1594.590 ;
        RECT 866.270 1594.530 869.170 1594.590 ;
        RECT 1046.270 1594.530 1049.170 1594.590 ;
        RECT 1226.270 1594.530 1229.170 1594.590 ;
        RECT 1406.270 1594.530 1409.170 1594.590 ;
        RECT 1586.270 1594.530 1589.170 1594.590 ;
        RECT 1766.270 1594.530 1769.170 1594.590 ;
        RECT 1946.270 1594.530 1949.170 1594.590 ;
        RECT 2126.270 1594.530 2129.170 1594.590 ;
        RECT 2306.270 1594.530 2309.170 1594.590 ;
        RECT 2486.270 1594.530 2489.170 1594.590 ;
        RECT 2666.270 1594.530 2669.170 1594.590 ;
        RECT 2846.270 1594.530 2849.170 1594.590 ;
        RECT 2958.850 1594.530 2961.750 1594.590 ;
        RECT -42.130 1591.630 2961.750 1594.530 ;
        RECT -42.130 1591.570 -39.230 1591.630 ;
        RECT 146.270 1591.570 149.170 1591.630 ;
        RECT 326.270 1591.570 329.170 1591.630 ;
        RECT 506.270 1591.570 509.170 1591.630 ;
        RECT 686.270 1591.570 689.170 1591.630 ;
        RECT 866.270 1591.570 869.170 1591.630 ;
        RECT 1046.270 1591.570 1049.170 1591.630 ;
        RECT 1226.270 1591.570 1229.170 1591.630 ;
        RECT 1406.270 1591.570 1409.170 1591.630 ;
        RECT 1586.270 1591.570 1589.170 1591.630 ;
        RECT 1766.270 1591.570 1769.170 1591.630 ;
        RECT 1946.270 1591.570 1949.170 1591.630 ;
        RECT 2126.270 1591.570 2129.170 1591.630 ;
        RECT 2306.270 1591.570 2309.170 1591.630 ;
        RECT 2486.270 1591.570 2489.170 1591.630 ;
        RECT 2666.270 1591.570 2669.170 1591.630 ;
        RECT 2846.270 1591.570 2849.170 1591.630 ;
        RECT 2958.850 1591.570 2961.750 1591.630 ;
        RECT -42.130 1414.530 -39.230 1414.590 ;
        RECT 146.270 1414.530 149.170 1414.590 ;
        RECT 326.270 1414.530 329.170 1414.590 ;
        RECT 506.270 1414.530 509.170 1414.590 ;
        RECT 686.270 1414.530 689.170 1414.590 ;
        RECT 866.270 1414.530 869.170 1414.590 ;
        RECT 1046.270 1414.530 1049.170 1414.590 ;
        RECT 1226.270 1414.530 1229.170 1414.590 ;
        RECT 1406.270 1414.530 1409.170 1414.590 ;
        RECT 1586.270 1414.530 1589.170 1414.590 ;
        RECT 1766.270 1414.530 1769.170 1414.590 ;
        RECT 1946.270 1414.530 1949.170 1414.590 ;
        RECT 2126.270 1414.530 2129.170 1414.590 ;
        RECT 2306.270 1414.530 2309.170 1414.590 ;
        RECT 2486.270 1414.530 2489.170 1414.590 ;
        RECT 2666.270 1414.530 2669.170 1414.590 ;
        RECT 2846.270 1414.530 2849.170 1414.590 ;
        RECT 2958.850 1414.530 2961.750 1414.590 ;
        RECT -42.130 1411.630 2961.750 1414.530 ;
        RECT -42.130 1411.570 -39.230 1411.630 ;
        RECT 146.270 1411.570 149.170 1411.630 ;
        RECT 326.270 1411.570 329.170 1411.630 ;
        RECT 506.270 1411.570 509.170 1411.630 ;
        RECT 686.270 1411.570 689.170 1411.630 ;
        RECT 866.270 1411.570 869.170 1411.630 ;
        RECT 1046.270 1411.570 1049.170 1411.630 ;
        RECT 1226.270 1411.570 1229.170 1411.630 ;
        RECT 1406.270 1411.570 1409.170 1411.630 ;
        RECT 1586.270 1411.570 1589.170 1411.630 ;
        RECT 1766.270 1411.570 1769.170 1411.630 ;
        RECT 1946.270 1411.570 1949.170 1411.630 ;
        RECT 2126.270 1411.570 2129.170 1411.630 ;
        RECT 2306.270 1411.570 2309.170 1411.630 ;
        RECT 2486.270 1411.570 2489.170 1411.630 ;
        RECT 2666.270 1411.570 2669.170 1411.630 ;
        RECT 2846.270 1411.570 2849.170 1411.630 ;
        RECT 2958.850 1411.570 2961.750 1411.630 ;
        RECT -42.130 1234.530 -39.230 1234.590 ;
        RECT 146.270 1234.530 149.170 1234.590 ;
        RECT 326.270 1234.530 329.170 1234.590 ;
        RECT 506.270 1234.530 509.170 1234.590 ;
        RECT 686.270 1234.530 689.170 1234.590 ;
        RECT 866.270 1234.530 869.170 1234.590 ;
        RECT 1046.270 1234.530 1049.170 1234.590 ;
        RECT 1226.270 1234.530 1229.170 1234.590 ;
        RECT 1406.270 1234.530 1409.170 1234.590 ;
        RECT 1586.270 1234.530 1589.170 1234.590 ;
        RECT 1766.270 1234.530 1769.170 1234.590 ;
        RECT 1946.270 1234.530 1949.170 1234.590 ;
        RECT 2126.270 1234.530 2129.170 1234.590 ;
        RECT 2306.270 1234.530 2309.170 1234.590 ;
        RECT 2486.270 1234.530 2489.170 1234.590 ;
        RECT 2666.270 1234.530 2669.170 1234.590 ;
        RECT 2846.270 1234.530 2849.170 1234.590 ;
        RECT 2958.850 1234.530 2961.750 1234.590 ;
        RECT -42.130 1231.630 2961.750 1234.530 ;
        RECT -42.130 1231.570 -39.230 1231.630 ;
        RECT 146.270 1231.570 149.170 1231.630 ;
        RECT 326.270 1231.570 329.170 1231.630 ;
        RECT 506.270 1231.570 509.170 1231.630 ;
        RECT 686.270 1231.570 689.170 1231.630 ;
        RECT 866.270 1231.570 869.170 1231.630 ;
        RECT 1046.270 1231.570 1049.170 1231.630 ;
        RECT 1226.270 1231.570 1229.170 1231.630 ;
        RECT 1406.270 1231.570 1409.170 1231.630 ;
        RECT 1586.270 1231.570 1589.170 1231.630 ;
        RECT 1766.270 1231.570 1769.170 1231.630 ;
        RECT 1946.270 1231.570 1949.170 1231.630 ;
        RECT 2126.270 1231.570 2129.170 1231.630 ;
        RECT 2306.270 1231.570 2309.170 1231.630 ;
        RECT 2486.270 1231.570 2489.170 1231.630 ;
        RECT 2666.270 1231.570 2669.170 1231.630 ;
        RECT 2846.270 1231.570 2849.170 1231.630 ;
        RECT 2958.850 1231.570 2961.750 1231.630 ;
        RECT -42.130 1054.530 -39.230 1054.590 ;
        RECT 146.270 1054.530 149.170 1054.590 ;
        RECT 326.270 1054.530 329.170 1054.590 ;
        RECT 506.270 1054.530 509.170 1054.590 ;
        RECT 686.270 1054.530 689.170 1054.590 ;
        RECT 866.270 1054.530 869.170 1054.590 ;
        RECT 1046.270 1054.530 1049.170 1054.590 ;
        RECT 1226.270 1054.530 1229.170 1054.590 ;
        RECT 1406.270 1054.530 1409.170 1054.590 ;
        RECT 1586.270 1054.530 1589.170 1054.590 ;
        RECT 1766.270 1054.530 1769.170 1054.590 ;
        RECT 1946.270 1054.530 1949.170 1054.590 ;
        RECT 2126.270 1054.530 2129.170 1054.590 ;
        RECT 2306.270 1054.530 2309.170 1054.590 ;
        RECT 2486.270 1054.530 2489.170 1054.590 ;
        RECT 2666.270 1054.530 2669.170 1054.590 ;
        RECT 2846.270 1054.530 2849.170 1054.590 ;
        RECT 2958.850 1054.530 2961.750 1054.590 ;
        RECT -42.130 1051.630 2961.750 1054.530 ;
        RECT -42.130 1051.570 -39.230 1051.630 ;
        RECT 146.270 1051.570 149.170 1051.630 ;
        RECT 326.270 1051.570 329.170 1051.630 ;
        RECT 506.270 1051.570 509.170 1051.630 ;
        RECT 686.270 1051.570 689.170 1051.630 ;
        RECT 866.270 1051.570 869.170 1051.630 ;
        RECT 1046.270 1051.570 1049.170 1051.630 ;
        RECT 1226.270 1051.570 1229.170 1051.630 ;
        RECT 1406.270 1051.570 1409.170 1051.630 ;
        RECT 1586.270 1051.570 1589.170 1051.630 ;
        RECT 1766.270 1051.570 1769.170 1051.630 ;
        RECT 1946.270 1051.570 1949.170 1051.630 ;
        RECT 2126.270 1051.570 2129.170 1051.630 ;
        RECT 2306.270 1051.570 2309.170 1051.630 ;
        RECT 2486.270 1051.570 2489.170 1051.630 ;
        RECT 2666.270 1051.570 2669.170 1051.630 ;
        RECT 2846.270 1051.570 2849.170 1051.630 ;
        RECT 2958.850 1051.570 2961.750 1051.630 ;
        RECT -42.130 874.530 -39.230 874.590 ;
        RECT 146.270 874.530 149.170 874.590 ;
        RECT 326.270 874.530 329.170 874.590 ;
        RECT 506.270 874.530 509.170 874.590 ;
        RECT 686.270 874.530 689.170 874.590 ;
        RECT 866.270 874.530 869.170 874.590 ;
        RECT 1046.270 874.530 1049.170 874.590 ;
        RECT 1226.270 874.530 1229.170 874.590 ;
        RECT 1406.270 874.530 1409.170 874.590 ;
        RECT 1586.270 874.530 1589.170 874.590 ;
        RECT 1766.270 874.530 1769.170 874.590 ;
        RECT 1946.270 874.530 1949.170 874.590 ;
        RECT 2126.270 874.530 2129.170 874.590 ;
        RECT 2306.270 874.530 2309.170 874.590 ;
        RECT 2486.270 874.530 2489.170 874.590 ;
        RECT 2666.270 874.530 2669.170 874.590 ;
        RECT 2846.270 874.530 2849.170 874.590 ;
        RECT 2958.850 874.530 2961.750 874.590 ;
        RECT -42.130 871.630 2961.750 874.530 ;
        RECT -42.130 871.570 -39.230 871.630 ;
        RECT 146.270 871.570 149.170 871.630 ;
        RECT 326.270 871.570 329.170 871.630 ;
        RECT 506.270 871.570 509.170 871.630 ;
        RECT 686.270 871.570 689.170 871.630 ;
        RECT 866.270 871.570 869.170 871.630 ;
        RECT 1046.270 871.570 1049.170 871.630 ;
        RECT 1226.270 871.570 1229.170 871.630 ;
        RECT 1406.270 871.570 1409.170 871.630 ;
        RECT 1586.270 871.570 1589.170 871.630 ;
        RECT 1766.270 871.570 1769.170 871.630 ;
        RECT 1946.270 871.570 1949.170 871.630 ;
        RECT 2126.270 871.570 2129.170 871.630 ;
        RECT 2306.270 871.570 2309.170 871.630 ;
        RECT 2486.270 871.570 2489.170 871.630 ;
        RECT 2666.270 871.570 2669.170 871.630 ;
        RECT 2846.270 871.570 2849.170 871.630 ;
        RECT 2958.850 871.570 2961.750 871.630 ;
        RECT -42.130 694.530 -39.230 694.590 ;
        RECT 146.270 694.530 149.170 694.590 ;
        RECT 326.270 694.530 329.170 694.590 ;
        RECT 506.270 694.530 509.170 694.590 ;
        RECT 686.270 694.530 689.170 694.590 ;
        RECT 866.270 694.530 869.170 694.590 ;
        RECT 1046.270 694.530 1049.170 694.590 ;
        RECT 1226.270 694.530 1229.170 694.590 ;
        RECT 1406.270 694.530 1409.170 694.590 ;
        RECT 1586.270 694.530 1589.170 694.590 ;
        RECT 1766.270 694.530 1769.170 694.590 ;
        RECT 1946.270 694.530 1949.170 694.590 ;
        RECT 2126.270 694.530 2129.170 694.590 ;
        RECT 2306.270 694.530 2309.170 694.590 ;
        RECT 2486.270 694.530 2489.170 694.590 ;
        RECT 2666.270 694.530 2669.170 694.590 ;
        RECT 2846.270 694.530 2849.170 694.590 ;
        RECT 2958.850 694.530 2961.750 694.590 ;
        RECT -42.130 691.630 2961.750 694.530 ;
        RECT -42.130 691.570 -39.230 691.630 ;
        RECT 146.270 691.570 149.170 691.630 ;
        RECT 326.270 691.570 329.170 691.630 ;
        RECT 506.270 691.570 509.170 691.630 ;
        RECT 686.270 691.570 689.170 691.630 ;
        RECT 866.270 691.570 869.170 691.630 ;
        RECT 1046.270 691.570 1049.170 691.630 ;
        RECT 1226.270 691.570 1229.170 691.630 ;
        RECT 1406.270 691.570 1409.170 691.630 ;
        RECT 1586.270 691.570 1589.170 691.630 ;
        RECT 1766.270 691.570 1769.170 691.630 ;
        RECT 1946.270 691.570 1949.170 691.630 ;
        RECT 2126.270 691.570 2129.170 691.630 ;
        RECT 2306.270 691.570 2309.170 691.630 ;
        RECT 2486.270 691.570 2489.170 691.630 ;
        RECT 2666.270 691.570 2669.170 691.630 ;
        RECT 2846.270 691.570 2849.170 691.630 ;
        RECT 2958.850 691.570 2961.750 691.630 ;
        RECT -42.130 514.530 -39.230 514.590 ;
        RECT 146.270 514.530 149.170 514.590 ;
        RECT 326.270 514.530 329.170 514.590 ;
        RECT 506.270 514.530 509.170 514.590 ;
        RECT 686.270 514.530 689.170 514.590 ;
        RECT 866.270 514.530 869.170 514.590 ;
        RECT 1046.270 514.530 1049.170 514.590 ;
        RECT 1226.270 514.530 1229.170 514.590 ;
        RECT 1406.270 514.530 1409.170 514.590 ;
        RECT 1586.270 514.530 1589.170 514.590 ;
        RECT 1766.270 514.530 1769.170 514.590 ;
        RECT 1946.270 514.530 1949.170 514.590 ;
        RECT 2126.270 514.530 2129.170 514.590 ;
        RECT 2306.270 514.530 2309.170 514.590 ;
        RECT 2486.270 514.530 2489.170 514.590 ;
        RECT 2666.270 514.530 2669.170 514.590 ;
        RECT 2846.270 514.530 2849.170 514.590 ;
        RECT 2958.850 514.530 2961.750 514.590 ;
        RECT -42.130 511.630 2961.750 514.530 ;
        RECT -42.130 511.570 -39.230 511.630 ;
        RECT 146.270 511.570 149.170 511.630 ;
        RECT 326.270 511.570 329.170 511.630 ;
        RECT 506.270 511.570 509.170 511.630 ;
        RECT 686.270 511.570 689.170 511.630 ;
        RECT 866.270 511.570 869.170 511.630 ;
        RECT 1046.270 511.570 1049.170 511.630 ;
        RECT 1226.270 511.570 1229.170 511.630 ;
        RECT 1406.270 511.570 1409.170 511.630 ;
        RECT 1586.270 511.570 1589.170 511.630 ;
        RECT 1766.270 511.570 1769.170 511.630 ;
        RECT 1946.270 511.570 1949.170 511.630 ;
        RECT 2126.270 511.570 2129.170 511.630 ;
        RECT 2306.270 511.570 2309.170 511.630 ;
        RECT 2486.270 511.570 2489.170 511.630 ;
        RECT 2666.270 511.570 2669.170 511.630 ;
        RECT 2846.270 511.570 2849.170 511.630 ;
        RECT 2958.850 511.570 2961.750 511.630 ;
        RECT -42.130 334.530 -39.230 334.590 ;
        RECT 146.270 334.530 149.170 334.590 ;
        RECT 326.270 334.530 329.170 334.590 ;
        RECT 506.270 334.530 509.170 334.590 ;
        RECT 686.270 334.530 689.170 334.590 ;
        RECT 866.270 334.530 869.170 334.590 ;
        RECT 1046.270 334.530 1049.170 334.590 ;
        RECT 1226.270 334.530 1229.170 334.590 ;
        RECT 1406.270 334.530 1409.170 334.590 ;
        RECT 1586.270 334.530 1589.170 334.590 ;
        RECT 1766.270 334.530 1769.170 334.590 ;
        RECT 1946.270 334.530 1949.170 334.590 ;
        RECT 2126.270 334.530 2129.170 334.590 ;
        RECT 2306.270 334.530 2309.170 334.590 ;
        RECT 2486.270 334.530 2489.170 334.590 ;
        RECT 2666.270 334.530 2669.170 334.590 ;
        RECT 2846.270 334.530 2849.170 334.590 ;
        RECT 2958.850 334.530 2961.750 334.590 ;
        RECT -42.130 331.630 2961.750 334.530 ;
        RECT -42.130 331.570 -39.230 331.630 ;
        RECT 146.270 331.570 149.170 331.630 ;
        RECT 326.270 331.570 329.170 331.630 ;
        RECT 506.270 331.570 509.170 331.630 ;
        RECT 686.270 331.570 689.170 331.630 ;
        RECT 866.270 331.570 869.170 331.630 ;
        RECT 1046.270 331.570 1049.170 331.630 ;
        RECT 1226.270 331.570 1229.170 331.630 ;
        RECT 1406.270 331.570 1409.170 331.630 ;
        RECT 1586.270 331.570 1589.170 331.630 ;
        RECT 1766.270 331.570 1769.170 331.630 ;
        RECT 1946.270 331.570 1949.170 331.630 ;
        RECT 2126.270 331.570 2129.170 331.630 ;
        RECT 2306.270 331.570 2309.170 331.630 ;
        RECT 2486.270 331.570 2489.170 331.630 ;
        RECT 2666.270 331.570 2669.170 331.630 ;
        RECT 2846.270 331.570 2849.170 331.630 ;
        RECT 2958.850 331.570 2961.750 331.630 ;
        RECT -42.130 154.530 -39.230 154.590 ;
        RECT 146.270 154.530 149.170 154.590 ;
        RECT 326.270 154.530 329.170 154.590 ;
        RECT 506.270 154.530 509.170 154.590 ;
        RECT 686.270 154.530 689.170 154.590 ;
        RECT 866.270 154.530 869.170 154.590 ;
        RECT 1046.270 154.530 1049.170 154.590 ;
        RECT 1226.270 154.530 1229.170 154.590 ;
        RECT 1406.270 154.530 1409.170 154.590 ;
        RECT 1586.270 154.530 1589.170 154.590 ;
        RECT 1766.270 154.530 1769.170 154.590 ;
        RECT 1946.270 154.530 1949.170 154.590 ;
        RECT 2126.270 154.530 2129.170 154.590 ;
        RECT 2306.270 154.530 2309.170 154.590 ;
        RECT 2486.270 154.530 2489.170 154.590 ;
        RECT 2666.270 154.530 2669.170 154.590 ;
        RECT 2846.270 154.530 2849.170 154.590 ;
        RECT 2958.850 154.530 2961.750 154.590 ;
        RECT -42.130 151.630 2961.750 154.530 ;
        RECT -42.130 151.570 -39.230 151.630 ;
        RECT 146.270 151.570 149.170 151.630 ;
        RECT 326.270 151.570 329.170 151.630 ;
        RECT 506.270 151.570 509.170 151.630 ;
        RECT 686.270 151.570 689.170 151.630 ;
        RECT 866.270 151.570 869.170 151.630 ;
        RECT 1046.270 151.570 1049.170 151.630 ;
        RECT 1226.270 151.570 1229.170 151.630 ;
        RECT 1406.270 151.570 1409.170 151.630 ;
        RECT 1586.270 151.570 1589.170 151.630 ;
        RECT 1766.270 151.570 1769.170 151.630 ;
        RECT 1946.270 151.570 1949.170 151.630 ;
        RECT 2126.270 151.570 2129.170 151.630 ;
        RECT 2306.270 151.570 2309.170 151.630 ;
        RECT 2486.270 151.570 2489.170 151.630 ;
        RECT 2666.270 151.570 2669.170 151.630 ;
        RECT 2846.270 151.570 2849.170 151.630 ;
        RECT 2958.850 151.570 2961.750 151.630 ;
        RECT -42.130 -33.870 -39.230 -33.810 ;
        RECT 146.270 -33.870 149.170 -33.810 ;
        RECT 326.270 -33.870 329.170 -33.810 ;
        RECT 506.270 -33.870 509.170 -33.810 ;
        RECT 686.270 -33.870 689.170 -33.810 ;
        RECT 866.270 -33.870 869.170 -33.810 ;
        RECT 1046.270 -33.870 1049.170 -33.810 ;
        RECT 1226.270 -33.870 1229.170 -33.810 ;
        RECT 1406.270 -33.870 1409.170 -33.810 ;
        RECT 1586.270 -33.870 1589.170 -33.810 ;
        RECT 1766.270 -33.870 1769.170 -33.810 ;
        RECT 1946.270 -33.870 1949.170 -33.810 ;
        RECT 2126.270 -33.870 2129.170 -33.810 ;
        RECT 2306.270 -33.870 2309.170 -33.810 ;
        RECT 2486.270 -33.870 2489.170 -33.810 ;
        RECT 2666.270 -33.870 2669.170 -33.810 ;
        RECT 2846.270 -33.870 2849.170 -33.810 ;
        RECT 2958.850 -33.870 2961.750 -33.810 ;
        RECT -42.130 -36.770 2961.750 -33.870 ;
        RECT -42.130 -36.830 -39.230 -36.770 ;
        RECT 146.270 -36.830 149.170 -36.770 ;
        RECT 326.270 -36.830 329.170 -36.770 ;
        RECT 506.270 -36.830 509.170 -36.770 ;
        RECT 686.270 -36.830 689.170 -36.770 ;
        RECT 866.270 -36.830 869.170 -36.770 ;
        RECT 1046.270 -36.830 1049.170 -36.770 ;
        RECT 1226.270 -36.830 1229.170 -36.770 ;
        RECT 1406.270 -36.830 1409.170 -36.770 ;
        RECT 1586.270 -36.830 1589.170 -36.770 ;
        RECT 1766.270 -36.830 1769.170 -36.770 ;
        RECT 1946.270 -36.830 1949.170 -36.770 ;
        RECT 2126.270 -36.830 2129.170 -36.770 ;
        RECT 2306.270 -36.830 2309.170 -36.770 ;
        RECT 2486.270 -36.830 2489.170 -36.770 ;
        RECT 2666.270 -36.830 2669.170 -36.770 ;
        RECT 2846.270 -36.830 2849.170 -36.770 ;
        RECT 2958.850 -36.830 2961.750 -36.770 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1156.520 1710.795 1795.460 2336.565 ;
      LAYER met1 ;
        RECT 1156.520 1710.640 1795.460 2336.720 ;
      LAYER met2 ;
        RECT 1168.110 2345.720 1196.810 2346.000 ;
        RECT 1197.650 2345.720 1289.270 2346.000 ;
        RECT 1290.110 2345.720 1382.190 2346.000 ;
        RECT 1383.030 2345.720 1475.110 2346.000 ;
        RECT 1475.950 2345.720 1568.030 2346.000 ;
        RECT 1568.870 2345.720 1660.950 2346.000 ;
        RECT 1661.790 2345.720 1753.870 2346.000 ;
        RECT 1754.710 2345.720 1788.010 2346.000 ;
        RECT 1168.110 1704.280 1788.010 2345.720 ;
        RECT 1168.110 1704.000 1191.290 1704.280 ;
        RECT 1192.130 1704.000 1272.250 1704.280 ;
        RECT 1273.090 1704.000 1353.670 1704.280 ;
        RECT 1354.510 1704.000 1434.630 1704.280 ;
        RECT 1435.470 1704.000 1516.050 1704.280 ;
        RECT 1516.890 1704.000 1597.470 1704.280 ;
        RECT 1598.310 1704.000 1678.430 1704.280 ;
        RECT 1679.270 1704.000 1759.850 1704.280 ;
        RECT 1760.690 1704.000 1788.010 1704.280 ;
      LAYER met3 ;
        RECT 1155.000 2314.400 1797.000 2336.645 ;
        RECT 1155.000 2313.000 1796.600 2314.400 ;
        RECT 1155.000 2242.320 1797.000 2313.000 ;
        RECT 1155.400 2240.920 1796.600 2242.320 ;
        RECT 1155.000 2170.240 1797.000 2240.920 ;
        RECT 1155.000 2168.840 1796.600 2170.240 ;
        RECT 1155.000 2098.160 1797.000 2168.840 ;
        RECT 1155.000 2096.760 1796.600 2098.160 ;
        RECT 1155.000 2025.400 1797.000 2096.760 ;
        RECT 1155.400 2024.000 1796.600 2025.400 ;
        RECT 1155.000 1953.320 1797.000 2024.000 ;
        RECT 1155.000 1951.920 1796.600 1953.320 ;
        RECT 1155.000 1881.240 1797.000 1951.920 ;
        RECT 1155.000 1879.840 1796.600 1881.240 ;
        RECT 1155.000 1809.160 1797.000 1879.840 ;
        RECT 1155.400 1807.760 1796.600 1809.160 ;
        RECT 1155.000 1737.080 1797.000 1807.760 ;
        RECT 1155.000 1735.680 1796.600 1737.080 ;
        RECT 1155.000 1710.715 1797.000 1735.680 ;
      LAYER met4 ;
        RECT 1169.720 1710.640 1171.320 2336.720 ;
        RECT 1259.720 1710.640 1261.320 2336.720 ;
      LAYER met4 ;
        RECT 1349.720 1710.640 1354.070 2336.720 ;
        RECT 1356.970 1710.640 1371.470 2336.720 ;
        RECT 1374.370 1710.640 1388.870 2336.720 ;
        RECT 1391.770 1710.640 1406.270 2336.720 ;
        RECT 1409.170 1710.640 1444.070 2336.720 ;
        RECT 1446.970 1710.640 1461.470 2336.720 ;
        RECT 1464.370 1710.640 1478.870 2336.720 ;
        RECT 1481.770 1710.640 1496.270 2336.720 ;
        RECT 1499.170 1710.640 1534.070 2336.720 ;
        RECT 1536.970 1710.640 1551.470 2336.720 ;
        RECT 1554.370 1710.640 1568.870 2336.720 ;
        RECT 1571.770 1710.640 1586.270 2336.720 ;
        RECT 1589.170 1710.640 1624.070 2336.720 ;
        RECT 1626.970 1710.640 1641.470 2336.720 ;
        RECT 1644.370 1710.640 1658.870 2336.720 ;
        RECT 1661.770 1710.640 1676.270 2336.720 ;
        RECT 1679.170 1710.640 1714.070 2336.720 ;
        RECT 1716.970 1710.640 1722.945 2336.720 ;
  END
END user_project_wrapper
END LIBRARY

