VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rapcore
  CLASS BLOCK ;
  FOREIGN rapcore ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 650.000 ;
  PIN BUFFER_DTR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 646.000 36.080 650.000 36.680 ;
    END
  END BUFFER_DTR
  PIN CHARGEPUMP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 646.000 46.370 650.000 ;
    END
  END CHARGEPUMP
  PIN CIPO
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 646.000 108.160 650.000 108.760 ;
    END
  END CIPO
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 646.000 180.240 650.000 180.840 ;
    END
  END CLK
  PIN COPI
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END COPI
  PIN CS
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END CS
  PIN DIRINPUT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.550 646.000 138.830 650.000 ;
    END
  END DIRINPUT
  PIN DIROUTPUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 646.000 252.320 650.000 252.920 ;
    END
  END DIROUTPUT
  PIN ENC_A
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END ENC_A
  PIN ENC_B
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END ENC_B
  PIN HALT
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END HALT
  PIN MOVE_DONE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END MOVE_DONE
  PIN PHASE_A1
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 646.000 324.400 650.000 325.000 ;
    END
  END PHASE_A1
  PIN PHASE_A1_H
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.470 646.000 231.750 650.000 ;
    END
  END PHASE_A1_H
  PIN PHASE_A2
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 646.000 397.160 650.000 397.760 ;
    END
  END PHASE_A2
  PIN PHASE_A2_H
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 324.390 646.000 324.670 650.000 ;
    END
  END PHASE_A2_H
  PIN PHASE_B1
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END PHASE_B1
  PIN PHASE_B1_H
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 646.000 469.240 650.000 469.840 ;
    END
  END PHASE_B1_H
  PIN PHASE_B2
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END PHASE_B2
  PIN PHASE_B2_H
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END PHASE_B2_H
  PIN SCK
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.310 646.000 417.590 650.000 ;
    END
  END SCK
  PIN STEPINPUT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 510.230 646.000 510.510 650.000 ;
    END
  END STEPINPUT
  PIN STEPOUTPUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END STEPOUTPUT
  PIN analog_cmp1
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.130 0.000 609.410 4.000 ;
    END
  END analog_cmp1
  PIN analog_cmp2
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 646.000 541.320 650.000 541.920 ;
    END
  END analog_cmp2
  PIN analog_out1
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 646.000 613.400 650.000 614.000 ;
    END
  END analog_out1
  PIN analog_out2
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.150 646.000 603.430 650.000 ;
    END
  END analog_out2
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.720 10.640 20.320 636.720 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 108.720 10.640 110.320 636.720 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 644.460 636.565 ;
      LAYER met1 ;
        RECT 5.520 10.640 644.460 636.720 ;
      LAYER met2 ;
        RECT 17.110 645.720 45.810 646.000 ;
        RECT 46.650 645.720 138.270 646.000 ;
        RECT 139.110 645.720 231.190 646.000 ;
        RECT 232.030 645.720 324.110 646.000 ;
        RECT 324.950 645.720 417.030 646.000 ;
        RECT 417.870 645.720 509.950 646.000 ;
        RECT 510.790 645.720 602.870 646.000 ;
        RECT 603.710 645.720 637.010 646.000 ;
        RECT 17.110 4.280 637.010 645.720 ;
        RECT 17.110 4.000 40.290 4.280 ;
        RECT 41.130 4.000 121.250 4.280 ;
        RECT 122.090 4.000 202.670 4.280 ;
        RECT 203.510 4.000 283.630 4.280 ;
        RECT 284.470 4.000 365.050 4.280 ;
        RECT 365.890 4.000 446.470 4.280 ;
        RECT 447.310 4.000 527.430 4.280 ;
        RECT 528.270 4.000 608.850 4.280 ;
        RECT 609.690 4.000 637.010 4.280 ;
      LAYER met3 ;
        RECT 4.000 614.400 646.000 636.645 ;
        RECT 4.000 613.000 645.600 614.400 ;
        RECT 4.000 542.320 646.000 613.000 ;
        RECT 4.400 540.920 645.600 542.320 ;
        RECT 4.000 470.240 646.000 540.920 ;
        RECT 4.000 468.840 645.600 470.240 ;
        RECT 4.000 398.160 646.000 468.840 ;
        RECT 4.000 396.760 645.600 398.160 ;
        RECT 4.000 325.400 646.000 396.760 ;
        RECT 4.400 324.000 645.600 325.400 ;
        RECT 4.000 253.320 646.000 324.000 ;
        RECT 4.000 251.920 645.600 253.320 ;
        RECT 4.000 181.240 646.000 251.920 ;
        RECT 4.000 179.840 645.600 181.240 ;
        RECT 4.000 109.160 646.000 179.840 ;
        RECT 4.400 107.760 645.600 109.160 ;
        RECT 4.000 37.080 646.000 107.760 ;
        RECT 4.000 35.680 645.600 37.080 ;
        RECT 4.000 10.715 646.000 35.680 ;
      LAYER met4 ;
        RECT 198.720 10.640 571.945 636.720 ;
  END
END rapcore
END LIBRARY

